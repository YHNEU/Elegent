-- Version: v11.9 11.9.0.4
-- File used only for Simulation

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Top_AD is

    port( sys_clk  : in    std_logic;
          sys_rest : in    std_logic;
          sts      : in    std_logic;
          data_in  : in    std_logic_vector(11 downto 0);
          rx_uart  : in    std_logic;
          ce       : out   std_logic;
          cs       : out   std_logic;
          rc       : out   std_logic;
          addr     : out   std_logic_vector(3 downto 0);
          tx_uart  : out   std_logic
        );

end Top_AD;

architecture DEF_ARCH of Top_AD is 

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOIN_IB
    port( YIN : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_TRI
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOTRI_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_IN
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DLN0P1C1
    port( D   : in    std_logic := 'U';
          G   : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKIO
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port(Y : out std_logic); 
  end component;

  component VCC
    port(Y : out std_logic); 
  end component;

    signal send_over, \data_recive[0]\, \data_recive[1]\, 
        \data_recive[2]\, \data_recive[3]\, \data_recive[4]\, 
        \data_recive[5]\, \data_recive[6]\, \data_recive[7]\, 
        receive_over, \data_ad[0]\, \data_ad[1]\, \data_ad[2]\, 
        \data_ad[3]\, \data_ad[4]\, \data_ad[5]\, \data_ad[6]\, 
        \data_ad[7]\, \data_ad[8]\, \data_ad[9]\, \data_ad[10]\, 
        \data_ad[11]\, ad_over, addr_over, send_whole_over, 
        conver_top, vld_whole, ad_once_over, receive_on, 
        \data_all[0]\, \data_all[1]\, \data_all[2]\, 
        \data_all[3]\, \data_all[4]\, \data_all[5]\, 
        \data_all[6]\, \data_all[7]\, \data_all[8]\, 
        \data_all[9]\, \data_all[10]\, \data_all[11]\, 
        \data_all[12]\, \data_all[13]\, \data_all[14]\, 
        \data_all[15]\, \data_all[16]\, \data_all[17]\, 
        \data_all[18]\, \data_all[19]\, \data_all[20]\, 
        \data_all[21]\, \data_all[22]\, \data_all[23]\, 
        \data_all[24]\, \data_all[25]\, \data_all[26]\, 
        \data_all[27]\, \data_all[28]\, \data_all[29]\, 
        \data_all[30]\, \data_all[31]\, \data_all[32]\, 
        \data_all[33]\, \data_all[34]\, \data_all[35]\, 
        \data_all[36]\, \data_all[37]\, \data_all[38]\, 
        \data_all[39]\, \data_all[40]\, \data_all[41]\, 
        \data_all[42]\, \data_all[43]\, \data_all[44]\, 
        \data_all[45]\, \data_all[46]\, \data_all[47]\, 
        \data_all[48]\, \data_all[49]\, \data_all[50]\, 
        \data_all[51]\, \data_all[52]\, \data_all[53]\, 
        \data_all[54]\, \data_all[55]\, \data_all[56]\, 
        \data_all[57]\, \data_all[58]\, \data_all[59]\, 
        \data_all[60]\, \data_all[61]\, \data_all[62]\, 
        \data_all[63]\, \data_all[64]\, \data_all[65]\, 
        \data_all[66]\, \data_all[67]\, \data_all[68]\, 
        \data_all[69]\, \data_all[70]\, \data_all[71]\, 
        \data_all[72]\, \data_all[73]\, \data_all[74]\, 
        \data_all[75]\, \data_all[76]\, \data_all[77]\, 
        \data_all[78]\, \data_all[79]\, \data_all[80]\, 
        \data_all[81]\, \data_all[82]\, \data_all[83]\, 
        \data_all[84]\, \data_all[85]\, \data_all[86]\, 
        \data_all[87]\, \data_all[88]\, \data_all[89]\, 
        \data_all[90]\, \data_all[91]\, \data_all[92]\, 
        \data_all[93]\, \data_all[94]\, \data_all[95]\, 
        \data_all[96]\, \data_all[97]\, \data_all[98]\, 
        \data_all[99]\, \data_all[100]\, \data_all[101]\, 
        \data_all[102]\, \data_all[103]\, \data_all[104]\, 
        \data_all[105]\, \data_all[106]\, \data_all[107]\, 
        \data_all[108]\, \data_all[109]\, \data_all[110]\, 
        \data_all[111]\, \data_all[112]\, \data_all[113]\, 
        \data_all[114]\, \data_all[115]\, \data_all[116]\, 
        \data_all[117]\, \data_all[118]\, \data_all[119]\, 
        \data_all[120]\, \data_all[121]\, \data_all[122]\, 
        \data_all[123]\, \data_all[124]\, \data_all[125]\, 
        \data_all[126]\, \data_all[127]\, \data_all[128]\, 
        \data_all[129]\, \data_all[130]\, \data_all[131]\, 
        \data_all[132]\, \data_all[133]\, \data_all[134]\, 
        \data_all[135]\, \data_all[136]\, \data_all[137]\, 
        \data_all[138]\, \data_all[139]\, \data_all[140]\, 
        \data_all[141]\, \data_all[142]\, \data_all[143]\, 
        \data_all[144]\, \data_all[145]\, \data_all[146]\, 
        \data_all[147]\, \data_all[148]\, \data_all[149]\, 
        \data_all[150]\, \data_all[151]\, \data_all[152]\, 
        \data_all[153]\, \data_all[154]\, \data_all[155]\, 
        \data_all[156]\, \data_all[157]\, \data_all[158]\, 
        \data_all[159]\, \data_all[160]\, \data_all[161]\, 
        \data_all[162]\, \data_all[163]\, \data_all[164]\, 
        \data_all[165]\, \data_all[166]\, \data_all[167]\, 
        \data_all[168]\, \data_all[169]\, \data_all[170]\, 
        \data_all[171]\, \data_all[172]\, \data_all[173]\, 
        \data_all[174]\, \data_all[175]\, \data_all[176]\, 
        \data_all[177]\, \data_all[178]\, \data_all[179]\, 
        \data_all[180]\, \data_all[181]\, \data_all[182]\, 
        \data_all[183]\, \data_all[184]\, \data_all[185]\, 
        \data_all[186]\, \data_all[187]\, \data_all[188]\, 
        \data_all[189]\, \data_all[190]\, \data_all[191]\, 
        \data_all[192]\, \data_all[193]\, \data_all[194]\, 
        \data_all[195]\, \data_all[196]\, \data_all[197]\, 
        \data_all[198]\, \data_all[199]\, \data_all[200]\, 
        \data_all[201]\, \data_all[202]\, \data_all[203]\, 
        \data_all[204]\, \data_all[205]\, \data_all[206]\, 
        \data_all[207]\, \data_all[208]\, \data_all[209]\, 
        \data_all[210]\, \data_all[211]\, \data_all[212]\, 
        \data_all[213]\, \data_all[214]\, \data_all[215]\, 
        \data_all[216]\, \data_all[217]\, \data_all[218]\, 
        \data_all[219]\, \data_all[220]\, \data_all[221]\, 
        \data_all[222]\, \data_all[223]\, \data_all[224]\, 
        \data_all[225]\, \data_all[226]\, \data_all[227]\, 
        \data_all[228]\, \data_all[229]\, \data_all[230]\, 
        \data_all[231]\, \data_all[232]\, \data_all[233]\, 
        \data_all[234]\, \data_all[235]\, \data_all[236]\, 
        \data_all[237]\, \data_all[238]\, \data_all[239]\, 
        vld_send, \data_send[0]\, \data_send[1]\, \data_send[2]\, 
        \data_send[3]\, \data_send[4]\, \data_send[5]\, 
        \data_send[6]\, \data_send[7]\, sys_clk_c, sys_rest_c, 
        sts_c, \data_in_c[0]\, \data_in_c[1]\, \data_in_c[2]\, 
        \data_in_c[3]\, \data_in_c[4]\, \data_in_c[5]\, 
        \data_in_c[6]\, \data_in_c[7]\, \data_in_c[8]\, 
        \data_in_c[9]\, \data_in_c[10]\, \data_in_c[11]\, 
        rx_uart_c, ce_c, rc_c, \addr_c[0]\, \addr_c[1]\, 
        \addr_c[2]\, \addr_c[3]\, tx_uart_c, \U4.N_31\, 
        addr_over_i, \addr_c_0[0]\, \U2/cnt_24_0_net_1\, 
        \U2/cnt[10]_net_1\, \U2/cnt_0_sqmuxa_net_1\, 
        \U2/un1_tx_uart27_1_1\, \U2/tx_uart36\, \U2/tx_uart27\, 
        \U2/un1_tx_uart27_6\, \U2/un1_tx_uart27_4_2\, 
        \U2/un1_tx_uart27_5\, \U2/un1_tx_uart27_4\, 
        \U2/un1_tx_uart27_0\, \U2/un1_tx_uart27_4_1\, 
        \U2/un1_tx_uart27_1_0\, \U2/N_111\, \U2/N_114\, 
        \U2/N_112\, \U2/tx_uart34_1\, \U2/N_194\, 
        \U2/tx_uart_11_iv_7\, \U2/data_send_m[7]\, 
        \U2/tx_uart_11_iv_1\, \U2/tx_uart_11_iv_3\, 
        \U2/tx_uart_11_iv_6\, \U2/parity_check_6_sqmuxa\, 
        \U2/tx_uart_11_iv_2\, \U2/tx_uart_11_iv_5\, 
        \U2/parity_check_1_sqmuxa\, \U2/data_send_m[2]\, 
        \U2/parity_check_5_sqmuxa\, \U2/data_send_m[6]\, 
        \U2/parity_check_2_sqmuxa\, \U2/data_send_m[3]\, 
        \U2/parity_check_net_1\, \U2/tx_uart_11_iv_0\, 
        \U2/tx_uart37_8\, \U2/tx_uart37_7\, \U2/send_net_1\, 
        \U2/parity_check_10_iv_0_4\, \U2/N_121\, \U2/N_119\, 
        \U2/parity_check_10_iv_0_1\, \U2/parity_check_10_iv_0_3\, 
        \U2/N_68_i\, \U2/parity_check_3_sqmuxa\, \U2/N_120\, 
        \U2/parity_check_10_iv_0_2\, \U2/N_60_i\, 
        \U2/parity_check_8_sqmuxa\, \U2/N_116\, \U2/N_55_i\, 
        \U2/parity_check_7_sqmuxa\, \U2/N_118\, \U2/tx_uart38_1\, 
        \U2/tx_uart37_6\, \U2/cnt[7]_net_1\, \U2/cnt[5]_net_1\, 
        \U2/tx_uart33_0_a2_0_2\, \U2/N_163\, \U2/un1_cnt_3\, 
        \U2/N_165\, \U2/cnt[8]_net_1\, \U2/tx_uart35_0_a2_0_1\, 
        \U2/N_166\, \U2/N_124\, \U2/tx_uart35_0_a2_0_0\, 
        \U2/cnt[3]_net_1\, \U2/cnt[0]_net_1\, 
        \U2/un1_tx_uart27_3_0_a2_3_1\, 
        \U2/un1_tx_uart27_3_0_a2_3_0\, \U2/cnt[6]_net_1\, 
        \U2/cnt[1]_net_1\, \U2/tx_uart36_8\, \U2/tx_uart36_5\, 
        \U2/tx_uart36_7\, \U2/un1_cnt_1\, \U2/cnt[4]_net_1\, 
        \U2/tx_uart36_6\, \U2/N_177\, \U2/cnt[2]_net_1\, 
        \U2/cnt[11]_net_1\, \U2/cnt[9]_net_1\, 
        \U2/tx_uart27_0_a2_3\, \U2/N_154\, \U2/tx_uart27_0_a2_2\, 
        \U2/tx_uart27_0_a2_1\, \U2/N_176\, \U2/tx_uart37_1\, 
        \U2/tx_uart37_0\, \U2/tx_uart37_6_0\, \U2/tx_uart37_3\, 
        \U2/tx_uart38_10_4\, \U2/N_7\, \U2/tx_uart38_10_3\, 
        \U2/tx_uart38_10_1\, \U2/N_129\, \U2/tx_uart34_0_a2_2_2\, 
        \U2/un1_cnt_4\, \U2/un1_cnt_8\, \U2/un1_cnt_2\, 
        \U2/un1_cnt_5\, \U2/N_169\, \U2/un1_tx_uart27_4_tz\, 
        \U2/un1_cnt\, \U2/tx_uart38\, \U2/tx_uart38_10\, 
        \U2/tx_uart_11\, \U2/N_196\, \U2/N_125\, 
        \U2/un1_tx_uart27\, \U2/parity_check_10_iv\, \U2/N_192\, 
        \U2/N_172\, \U2/N_197\, \U2/N_171\, \U2/N_181\, 
        \U2/N_180\, \U2/cnt_n3_net_1\, \U2/cnt_c2_net_1\, 
        \U2/cnt_n4_net_1\, \U2/cnt_n4_tz_net_1\, 
        \U2/cnt_n6_net_1\, \U2/cnt_n6_tz_net_1\, 
        \U2/cnt_c4_net_1\, \U2/cnt_n7_net_1\, \U2/cnt_c6_net_1\, 
        \U2/cnt_n9_net_1\, \U2/cnt_c8_net_1\, \U2/cnt_n10_net_1\, 
        \U2/cnt_c9_net_1\, \U2/cnt_n8_net_1\, \U2/cnt_c7_net_1\, 
        \U2/cnt_n5_net_1\, \U2/cnt_n2_net_1\, \U2/un5_vld_send\, 
        \U2/idle_send_net_1\, \U2/N_168\, \U2/N_127\, \U2/N_174\, 
        \U2/N_126\, \U2/N_153\, \U2/cnt_n11_net_1\, \U2/N_152\, 
        \U2/cnt_n1_net_1\, \U2/cnt_n0_net_1\, 
        \U2/idle_send_0_sqmuxa\, \U2/idle_send_2_sqmuxa\, 
        \U2/N_198\, \U2/parity_check_0_sqmuxa\, \U2/N_59_i\, 
        \U2/N_178\, \U2/N_173\, \U2/N_131\, \U2/N_128\, 
        \U2/N_164\, \U2/tx_uart_11_sqmuxa\, \U3/cnt[1]_net_1\, 
        \U3/cnt[0]_net_1\, \U3/cnt[3]_net_1\, 
        \U3/DWACT_FINC_E[0]\, \U3/cnt[8]_net_1\, 
        \U3/DWACT_FINC_E[4]\, \U3/recive_i\, \U3/recive_net_1\, 
        \U3/m87_0\, \U3/m81_0\, \U3/m91_0\, \U3/m72_0\, 
        \U3/m85_0\, \U3/m83_0\, \U3/m79_4\, \U3/m79_2\, 
        \U3/cnt[5]_net_1\, \U3/m79_3\, \U3/cnt[10]_net_1\, 
        \U3/cnt[7]_net_1\, \U3/m36_4\, \U3/m36_1\, \U3/m36_3\, 
        \U3/m89_0\, \U3/m93_0\, \U3/m27_2\, \U3/m27_1\, 
        \U3/m22_2\, \U3/m22_0\, \U3/m22_1\, \U3/m53_3\, 
        \U3/m53_2\, \U3/m47_3\, \U3/m47_1\, \U3/m47_2\, 
        \U3/m70_5\, \U3/m70_4\, \U3/cnt[2]_net_1\, \U3/m11_3\, 
        \U3/m62_6\, \U3/m62_4\, \U3/m62_5\, \U3/cnt[6]_net_1\, 
        \U3/m106_7\, \U3/m106_6\, \U3/m106_5\, \U3/m106_0\, 
        \U3/cnt[4]_net_1\, \U3/cnt[9]_net_1\, \U3/cnt[11]_net_1\, 
        \U3/m11_9\, \U3/m11_2\, \U3/m11_6\, \U3/m11_8\, 
        \U3/m11_4\, \U3/m17_1\, \U3/m17_0\, \U3/m41_0\, 
        \U3/data_recive29\, \U3/N_30_0\, \U3/data_recive26\, 
        \U3/data_recive24\, \U3/N_125_mux\, \U3/data_recive30\, 
        \U3/N_110_mux\, \U3/N_120_mux\, \U3/N_39\, 
        \U3/data_recive31\, \U3/data_recive28\, 
        \U3/data_recive27\, \U3/data_recive23\, 
        \U3/data_recive25\, \U3/N_29\, \U3/un1_cnt\, \U3/un2_cnt\, 
        \U3/rx_down_net_1\, \U3/idle_recive_i_0\, 
        \U3/data_recive_12[0]\, \U3/data_recive_12[2]\, 
        \U3/data_recive_12[4]\, \U3/data_recive_12[5]\, 
        \U3/receive_over_0_sqmuxa\, \U3/data_recive_12[7]\, 
        \U3/data_recive_12[6]\, \U3/data_recive_12[3]\, 
        \U3/cnt_4[0]\, \U3/cnt_4[7]_net_1\, \U3/cnt_4[6]_net_1\, 
        \U3/cnt_4[5]_net_1\, \U3/cnt_4[11]_net_1\, 
        \U3/cnt_4[3]_net_1\, \U3/data_recive_12[1]\, 
        \U3/rx_down_1\, \U3/rx_fall2_net_1\, \U3/rx_fall1_net_1\, 
        \U3/rx_fall_net_1\, \U3/I_5\, \U3/I_7\, \U3/I_12\, 
        \U3/I_23\, \U3/I_26\, \U3/I_28\, \U3/N_2\, 
        \U3/DWACT_FINC_E[6]\, \U3/DWACT_FINC_E[2]\, 
        \U3/DWACT_FINC_E[5]\, \U3/N_3\, \U3/DWACT_FINC_E[3]\, 
        \U3/N_5\, \U3/N_6\, \U3/N_7\, \U3/DWACT_FINC_E[1]\, 
        \U3/N_8\, \U3/N_10\, \U4/N_20\, \U4/N_7_0\, 
        \U4/conver_ris2_i\, \U4/conver_ris2_net_1\, \U4/N_23\, 
        \U4/N_22\, \U4/N_10_0\, \U4/conver_ris_net_1\, 
        \U4/pr_state[0]_net_1\, \U4/addr_n1\, \U4/addr_n2\, 
        \U4/N_8_0\, \U4/addr_n3\, \U4/N_9_0\, \U4/N_11_0\, 
        \U4/pr_state[1]_net_1\, \U4/N_6_0\, 
        \U4/nx_state_RNO[0]_net_1\, \U4/nx_state_RNO_0[0]_net_1\, 
        \U4/N_27\, \U4/N_25\, \U4/nx_state_RNO[1]_net_1\, 
        \U4/N_24\, \U4/nx_state_RNO_0[1]_net_1\, 
        \U4/conver_ris_2\, \U4/conver_ris3_i_0\, 
        \U4/conver_ris1_net_1\, \U4/nx_state[0]_net_1\, \GND\, 
        \U4/nx_state[1]_net_1\, \U1/pr_state_0[7]_net_1\, 
        \U1/pr_state_RNICDI39[1]_net_1\, \U1/pr_state_0[5]_net_1\, 
        \U1/N_119\, \U1/N_841_0\, \U1/m103_i_o2_0_o2_0_net_1\, 
        \U1/N_817\, \U1/N_831_0\, 
        \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_0[63]_net_1\, 
        \U1/N_833_0\, \U1/N_826\, \U1/N_819\, \U1/N_839_0\, 
        \U1/N_818\, \U1/N_835_0\, \U1/m302_0_i_o2_0_net_1\, 
        \U1/N_844_0\, \U1/data_all_3_i_0_0_o2_1[190]_net_1\, 
        \U1/N_830_0\, \U1/N_820\, \U1/N_838_0\, 
        \U1/m146_i_0_o2_1\, \U1/N_832_0\, 
        \U1/m253_i_0_o2_0_net_1\, \U1/N_842_0\, 
        \U1/m79_0_i_i_o2_0_net_1\, \U1/N_836_0\, 
        \U1/m125_0_0_i_o2_0_net_1\, \U1/N_837_0\, \U1/N_829_0\, 
        \U1/N_840_0\, \U1/N_834_0\, \U1/N_821\, \U1/N_1091\, 
        \U1/pr_state_RNIV2MS[1]_net_1\, \U1/pr_state[2]_net_1\, 
        \U1/pr_state_0[2]\, \U1/N_852\, \U1/cnt_daly[7]_net_1\, 
        \U1/cnt_daly[8]_net_1\, \U1/N_850\, \U1/N_810\, 
        \U1/pr_state[7]_net_1\, \U1/N_2303\, 
        \U1/cnt_daly[6]_net_1\, \U1/N_849\, 
        \U1/cnt_daly[5]_net_1\, \U1/N_848\, 
        \U1/cnt_daly[3]_net_1\, \U1/cnt_daly[4]_net_1\, 
        \U1/N_846\, \U1/cnt_daly[0]_net_1\, 
        \U1/cnt_daly[1]_net_1\, \U1/cnt_daly[2]_net_1\, 
        \U1/un2_data_filter[10]\, \U1/data_filter[10]_net_1\, 
        \U1/N319\, \U1/N_37\, \U1/data_filter_4_i_0_0_0[10]\, 
        \U1/I79_un1_Y\, \U1/ADD_14x14_fast_I79_Y_0\, 
        \U1/I64_un1_Y\, \U1/N262\, \U1/N269\, \U1/N246\, 
        \U1/N243\, \U1/N242\, \U1/data_filter[5]_net_1\, 
        \U1/N189\, \U1/data_filter[4]_net_1\, \U1/OVER\, 
        \U1/DWACT_FDEC_E[0]\, \U1/data_all_3_0_i_0_0[116]\, 
        \U1/N_830\, \U1/data_all_3_i_0_0_0[100]\, \U1/N_829\, 
        \U1/data_all_3_i_0_0_0[102]\, 
        \U1/data_all_3_0_i_0_0[125]\, 
        \U1/data_all_3_i_0_0_0[104]\, 
        \U1/data_all_3_i_0_0_0[105]\, 
        \U1/data_all_3_i_0_0_0[106]\, 
        \U1/data_all_3_i_0_0_0[107]\, 
        \U1/data_all_3_i_0_0_0[108]\, 
        \U1/data_all_3_0_i_0_0[120]\, \U1/data_all_3_i_0_0_0[96]\, 
        \U1/data_all_3_i_0_0_0[97]\, \U1/data_all_3_i_0_0_0[98]\, 
        \U1/data_all_3_i_0_0_0[99]\, \U1/data_all_3_i_0_0_0[101]\, 
        \U1/data_all_3_0_i_0_0[112]\, 
        \U1/data_all_3_i_0_0_0[103]\, 
        \U1/data_all_3_0_i_0_0[114]\, 
        \U1/data_all_3_0_i_0_0[115]\, 
        \U1/data_all_3_0_i_0_0[117]\, 
        \U1/data_all_3_0_i_0_0[118]\, 
        \U1/data_all_3_0_i_0_0[119]\, 
        \U1/data_all_3_i_0_0_0[109]\, 
        \U1/data_all_3_0_i_0_0[121]\, 
        \U1/data_all_3_0_i_0_0[122]\, 
        \U1/data_all_3_0_i_0_0[123]\, 
        \U1/data_all_3_0_i_0_0[124]\, 
        \U1/data_all_3_0_i_0_0[113]\, \U1/m252_i_0_0\, 
        \U1/m249_i_0_0\, \U1/m246_i_0_0\, 
        \U1/data_all_3_0_0_i_0[80]\, \U1/data_all_3_0_i_0_0[93]\, 
        \U1/m212_0_i_0\, \U1/N_833\, \U1/m237_i_0_0\, 
        \U1/data_all_3_0_0_i_0[83]\, \U1/m243_i_0_0\, 
        \U1/data_all_3_0_0_i_0[86]\, \U1/m225_i_0_0\, 
        \U1/m231_i_0_0\, \U1/data_all_3_0_0_i_0[85]\, 
        \U1/m228_i_0_0\, \U1/data_all_3_0_0_i_0[88]\, 
        \U1/m234_i_0_0\, \U1/data_all_3_0_i_0_0[185]\, \U1/N_844\, 
        \U1/data_all_3_0_i_0_0[178]\, 
        \U1/data_all_3_0_i_0_0[183]\, 
        \U1/data_all_3_0_i_0_0[184]\, \U1/data_all_3_0_i_0_0[61]\, 
        \U1/data_all_3_0_i_0_0[182]\, \U1/m205_0_i_0\, 
        \U1/m202_0_i_0\, \U1/N_841\, \U1/data_all_3_0_i_0_0[177]\, 
        \U1/data_all_3_0_i_0_0[141]\, \U1/data_all_3_0_0_i_0[60]\, 
        \U1/data_all_3_0_i_0_0[179]\, 
        \U1/data_all_3_0_i_0_0[133]\, 
        \U1/data_all_3_0_i_0_0[128]\, \U1/m199_0_i_0\, 
        \U1/data_all_3_0_i_0_0[134]\, \U1/data_all_3_0_0_i_0[48]\, 
        \U1/data_all_3_0_0_i_0[54]\, \U1/data_all_3_0_i_0_0[132]\, 
        \U1/data_all_3_0_i_0_0[129]\, 
        \U1/data_all_3_0_i_0_0[131]\, 
        \U1/data_all_3_0_i_0_0[188]\, 
        \U1/data_all_3_0_i_0_0[140]\, 
        \U1/data_all_3_0_i_0_0[137]\, 
        \U1/data_all_3_0_i_0_0[181]\, 
        \U1/data_all_3_0_i_0_0[139]\, 
        \U1/data_all_3_0_i_0_0[180]\, 
        \U1/data_all_3_0_i_0_0[176]\, 
        \U1/data_all_3_0_i_0_0[189]\, \U1/data_all_3_0_0_i_0[56]\, 
        \U1/data_all_3_0_0_i_0[52]\, \U1/data_all_3_0_0_i_0[53]\, 
        \U1/m147_0_0_i_0\, \U1/m141_0_i_0_0\, \U1/N_836\, 
        \U1/m150_i_0_0\, \U1/m82_1_i_i_0\, \U1/N_842\, 
        \U1/m92_1_i_0_0\, \U1/m95_1_i_0_0\, \U1/m138_0_i_0_0\, 
        \U1/m135_0_i_0_0\, \U1/m125_0_0_i_0\, \U1/m118_0_i_1_0\, 
        \U1/m286_i_0_0\, \U1/m103_0_i_0_0\, \U1/m112_1_i_0_0\, 
        \U1/m156_0_i_0_0\, \U1/m144_0_i_0_0\, \U1/m98_0_i_i_0\, 
        \U1/m79_0_i_i_0\, \U1/data_all_3_0_0_i_0[0]\, 
        \U1/m88_0_i_0_0\, \U1/m83_1_i_0_0\, \U1/m109_0_i_0_0\, 
        \U1/m106_0_i_0_0\, \U1/data_all_3_0_0_i_0[6]\, 
        \U1/data_all_3_0_0_i_0[13]\, \U1/m271_i_0_0\, \U1/N_832\, 
        \U1/m274_i_0_0\, \U1/m159_0_i_0_0\, \U1/m261_i_0_0\, 
        \U1/m289_i_0_0\, \U1/data_all_3_0_0_i_0[7]\, 
        \U1/m283_i_0_0\, \U1/data_all_3_0_0_i_0[8]\, \U1/N_835\, 
        \U1/data_all_3_0_0_i_0[12]\, \U1/data_all_3_0_0_i_0[4]\, 
        \U1/m280_i_0_0\, \U1/m298_i_0_0\, \U1/m292_i_0_0\, 
        \U1/m163_0_i_0_0\, \U1/m258_i_0_0\, \U1/m142_0_i_0\, 
        \U1/data_all_3_0_0_i_0[234]\, \U1/m136_i_0_0\, \U1/N_839\, 
        \U1/m130_0_i_0\, \U1/m121_0_0_i_0\, \U1/m145_i_0_0\, 
        \U1/m98_1_i_0\, \U1/m133_i_0_0\, \U1/m106_i_0_0\, 
        \U1/m139_0_i_0\, \U1/m124_0_i_0\, \U1/m89_i_0_0\, 
        \U1/m127_i_0_0\, \U1/m112_0_0_i_0\, 
        \U1/data_all_3_0_i_0_0[204]\, \U1/m82_0_i_0_0\, 
        \U1/m69_i_0_0\, \U1/data_all_3_i_0_0_0[224]\, 
        \U1/m118_0_i_0_0\, \U1/data_filter_4_i_0_0_0[8]\, 
        \U1/data_all_3_0_0_i_0[213]\, 
        \U1/data_all_3_0_i_0_0[210]\, 
        \U1/data_all_3_0_0_i_0[212]\, \U1/m57_0_i_0_0\, 
        \U1/data_all_3_0_0_i_0[214]\, 
        \U1/data_all_3_0_0_i_0[208]\, \U1/m64_1_i_0_0\, 
        \U1/data_all_3_0_i_0_0[218]\, 
        \U1/data_all_3_0_0_i_0[220]\, \U1/m188_i_0_0\, 
        \U1/m173_i_0_0\, \U1/N_838\, \U1/m153_i_0_0\, 
        \U1/m185_i_0_0\, \U1/m176_i_0_0\, \U1/m191_i_0_0\, 
        \U1/m156_i_0_0\, \U1/m161_i_0_0\, \U1/m179_i_0_0\, 
        \U1/m167_i_0_0\, \U1/m164_i_0_0\, \U1/m71_i_0_0\, 
        \U1/m170_i_0_0\, \U1/m182_i_0_0\, 
        \U1/data_filter_4_i_0_0_0[4]\, \U1/data_filter[6]_net_1\, 
        \U1/data_filter_4_i_0_0_0[11]\, 
        \U1/data_filter[13]_net_1\, \U1/pr_state[5]_net_1\, 
        \U1/data_filter[12]_net_1\, \U1/ADD_14x14_fast_I96_Y_0\, 
        \U1/data_filter[8]_net_1\, \U1/I_5_0\, \U1/I_9_0\, 
        \U1/m45_0_0_0\, \U1/data_filter[11]_net_1\, 
        \U1/ADD_14x14_fast_I77_Y_2\, \U1/N258\, \U1/N265\, 
        \U1/ADD_14x14_fast_I77_Y_1\, \U1/N231\, \U1/N234\, 
        \U1/ADD_14x14_fast_I77_Y_0\, \U1/N206\, \U1/m48_0_0_0\, 
        \U1/data_filter[9]_net_1\, \U1/m68_i_i_1\, \U1/N_870\, 
        \U1/N_866\, \U1/N_869\, \U1/m51_0_0_0\, \U1/m54_0_0_0\, 
        \U1/data_filter[7]_net_1\, \U1/m85_i_0_a3_1\, 
        \U1/pr_state[4]_net_1\, \U1/pr_state[3]_net_1\, 
        \U1/ADD_14x14_fast_I99_Y_0\, 
        \U1/ADD_14x14_fast_I77_un1_Y_0\, \U1/N239\, 
        \U1/ADD_14x14_fast_I76_Y_1\, \U1/N256\, \U1/N263\, 
        \U1/ADD_14x14_fast_I76_Y_0\, \U1/N229\, \U1/N232\, 
        \U1/N227\, \U1/I_7_0\, \U1/data_filter_4_i_0_0_0[3]\, 
        \U1/data_filter_4_i_0_0_0[2]\, 
        \U1/ADD_14x14_fast_I78_Y_1\, 
        \U1/ADD_14x14_fast_I78_un1_Y_0\, \U1/N275\, 
        \U1/ADD_14x14_fast_I78_Y_0\, \U1/N236\, \U1/N233\, 
        \U1/N238\, \U1/N235\, \U1/ADD_14x14_fast_I76_un1_Y_0\, 
        \U1/N264\, \U1/ADD_14x14_fast_I80_Y_0\, 
        \U1/ADD_14x14_fast_I80_un1_Y_0\, \U1/N237\, \U1/N268\, 
        \U1/N245\, \U1/N249\, \U1/N176\, \U1/m57_0_0_0\, 
        \U1/data_filter[3]_net_1\, \U1/m22_m4_0_a2_4\, 
        \U1/m22_m4_0_a2_2\, \U1/m22_m4_0_a2_3\, 
        \U1/cnt_daly[9]_net_1\, \U1/m77_i_0_0\, \U1/N_1084\, 
        \U1/N_878\, \U1/m61_0_i_a3_1_9\, \U1/m61_0_i_a3_1_1\, 
        \U1/m61_0_i_a3_1_0\, \U1/m61_0_i_a3_1_5\, 
        \U1/m61_0_i_a3_1_8\, \U1/m24_m4_e_2\, \U1/m61_0_i_a3_1_7\, 
        \U1/m61_0_i_a3_1_2\, \U1/pr_state[0]_net_1\, 
        \U1/cnt_daly[11]_net_1\, \U1/cnt_daly[12]_net_1\, 
        \U1/cnt_daly[10]_net_1\, \U1/m101_i_0_a3_0_0\, 
        \U1/m20_m6_0_a2_7\, \U1/m20_m6_0_a2_2\, 
        \U1/m20_m6_0_a2_1\, \U1/N_845\, \U1/m20_m6_0_a2_6\, 
        \U1/m20_m6_0_a2_4\, \U1/m24_m4_e_4\, \U1/m24_m4_e_3\, 
        \U1/m112_i_0_a3_0\, \U1/cnt_receive_over_net_1\, 
        \U1/m110_i_0_a3_1\, \U1/receive_flag_net_1\, 
        \U1/m107_e_3_net_1\, \U1/m107_e_2_net_1\, 
        \U1/m107_e_1_net_1\, \U1/N_840\, \U1/N_837\, \U1/N_831\, 
        \U1/m24_N_11_mux\, \U1/m22_N_11_mux\, \U1/m20_N_13_mux\, 
        \U1/N_765\, \U1/N_2253\, \U1/N_2254\, \U1/N_744\, 
        \U1/N_1809\, \U1/N_290\, \U1/N_315\, \U1/N_331\, 
        \U1/N_694\, \U1/N_372\, \U1/N_388\, \U1/N_401\, 
        \U1/N_417\, \U1/N_255\, \U1/N_239\, \U1/N_94\, \U1/N_100\, 
        \U1/N_187\, \U1/N_955\, \U1/N_956\, \U1/N_31\, \U1/N_245\, 
        \U1/N_139\, \U1/N_1780\, \U1/N_390\, \U1/N_403\, 
        \U1/N_419\, \U1/N_166\, \U1/N_56\, \U1/N_213\, \U1/N_217\, 
        \U1/N_227\, \U1/N_256\, \U1/N_860\, \U1/N_856\, 
        \U1/pr_state[6]_net_1\, \U1/N_796\, \U1/N_798\, 
        \U1/N_800\, \U1/N_802\, \U1/N_2299\, \U1/N_804\, 
        \U1/N_806\, \U1/N_808\, \U1/cnt[2]_net_1\, 
        \U1/cnt[0]_net_1\, \U1/cnt[1]_net_1\, \U1/N_871\, 
        \U1/N_857\, \U1/pr_state[1]_net_1\, \U1/N_1095\, 
        \U1/un2_data_filter[1]\, \U1/data_filter[1]_net_1\, 
        \U1/un2_data_filter[3]\, \U1/un2_data_filter[4]\, 
        \U1/N273\, \U1/un2_data_filter[5]\, \U1/N332\, 
        \U1/un2_data_filter[6]\, \U1/N329\, 
        \U1/un2_data_filter[7]\, \U1/N326\, 
        \U1/un2_data_filter[8]\, \U1/I68_un1_Y\, 
        \U1/un2_data_filter[9]\, \U1/N321\, 
        \U1/un2_data_filter[11]\, \U1/I62_un1_Y\, 
        \U1/un2_data_filter[2]\, \U1/data_filter[2]_net_1\, 
        \U1/N250\, \U1/N_854\, \U1/pr_state_RNO[0]_net_1\, 
        \U1/N_864\, \U1/N_865\, \U1/N_252\, \U1/N_41\, 
        \U1/N_1421\, \U1/N_45\, \U1/N_49\, \U1/N_1422\, \U1/N_43\, 
        \U1/N_48\, \U1/N_46_0\, \U1/N_49_0\, \U1/N_52_0\, 
        \U1/N_55_0\, \U1/N_58_0\, \U1/N_61_0\, \U1/N_906\, 
        \U1/N_905\, \U1/N_225\, \U1/N_909\, \U1/N_910\, 
        \U1/N_223\, \U1/N_911\, \U1/N_912\, \U1/N_221\, 
        \U1/N_219\, \U1/N_915\, \U1/N_916\, \U1/N_215\, 
        \U1/N_919\, \U1/N_920\, \U1/N_75\, \U1/N_77\, \U1/N_925\, 
        \U1/N_926\, \U1/N_2041\, \U1/N_2042\, \U1/N_85\, 
        \U1/N_206\, \U1/N_89\, \U1/N_203\, \U1/N_201\, \U1/N_93\, 
        \U1/N_96\, \U1/N_197\, \U1/data_filter[0]_net_1\, 
        \U1/N_101\, \U1/N_947\, \U1/N_948\, \U1/N_103\, 
        \U1/N_105\, \U1/N_107\, \U1/N_185\, \U1/N_957\, 
        \U1/N_958\, \U1/N_183\, \U1/N_959\, \U1/N_960\, 
        \U1/N_181\, \U1/N_179\, \U1/N_177\, \U1/N_175\, 
        \U1/N_173\, \U1/N_171\, \U1/N_971\, \U1/N_972\, 
        \U1/N_169\, \U1/N_167\, \U1/N_165\, \U1/N_163\, 
        \U1/N_2043\, \U1/N_981\, \U1/N_982\, \U1/N_160\, 
        \U1/N_30\, \U1/N_983\, \U1/N_984\, \U1/N_32\, \U1/N_985\, 
        \U1/N_986\, \U1/N_34\, \U1/N_1608\, \U1/N_1609\, 
        \U1/N_1611\, \U1/N_44\, \U1/N_46\, \U1/N_1612\, \U1/N_50\, 
        \U1/N_52\, \U1/N_54\, \U1/N_58\, \U1/N_60\, \U1/N_1613\, 
        \U1/N_1614\, \U1/N_1615\, \U1/N_170\, \U1/N_1017\, 
        \U1/N_1018\, \U1/N_174\, \U1/N_1019\, \U1/N_1020\, 
        \U1/N_178\, \U1/N_1021\, \U1/N_1022\, \U1/N_182\, 
        \U1/N_186\, \U1/N_190\, \U1/N_192\, \U1/N_1029\, 
        \U1/N_1030\, \U1/N_194\, \U1/N_1031\, \U1/N_1032\, 
        \U1/N_196\, \U1/N_199\, \U1/N_1035\, \U1/N_1036\, 
        \U1/N_202\, \U1/N_205\, \U1/N_208\, \U1/N_210\, 
        \U1/N_1043\, \U1/N_1044\, \U1/N_212\, \U1/N_216\, 
        \U1/N_1047\, \U1/N_1048\, \U1/N_220\, \U1/N_2073\, 
        \U1/N_1050\, \U1/N_224\, \U1/N_19\, \U1/N_97\, 
        \U1/N_1837\, \U1/N_87\, \U1/N_82\, \U1/N_1836\, \U1/N_78\, 
        \U1/N_73\, \U1/N_1835\, \U1/N_241\, \U1/N_1075\, 
        \U1/N_1076\, \U1/N_243\, \U1/N_1077\, \U1/N_1078\, 
        \U1/N_246\, \U1/N_248\, \U1/N_250\, \U1/N_253\, 
        \U1/N_1086\, \U1/N_1087\, \U1/N_258\, \U1/N_1096\, 
        \U1/N_1097\, \U1/N_261\, \U1/N_1098\, \U1/N_1099\, 
        \U1/N_264\, \U1/N_35\, \U1/N_39\, \U1/N_304\, \U1/N_53\, 
        \U1/N_415\, \U1/N_2079\, \U1/N_2080\, \U1/N_413\, 
        \U1/N_2081\, \U1/N_2082\, \U1/N_411\, \U1/N_409\, 
        \U1/N_407\, \U1/N_405\, \U1/N_399\, \U1/N_397\, 
        \U1/N_395\, \U1/N_393\, \U1/N_72\, \U1/N_386\, \U1/N_384\, 
        \U1/N_382\, \U1/N_380\, \U1/N_378\, \U1/N_376\, 
        \U1/N_374\, \U1/N_370\, \U1/N_368\, \U1/N_366\, 
        \U1/N_364\, \U1/N_362\, \U1/N_2131\, \U1/N_2132\, 
        \U1/N_360\, \U1/N_2133\, \U1/N_2134\, \U1/N_358\, 
        \U1/N_2135\, \U1/N_2136\, \U1/N_356\, \U1/N_680\, 
        \U1/N_2139\, \U1/N_2140\, \U1/N_686\, \U1/N_2141\, 
        \U1/N_2142\, \U1/N_688\, \U1/N_2143\, \U1/N_2144\, 
        \U1/N_690\, \U1/N_692\, \U1/N_2147\, \U1/N_2148\, 
        \U1/N_696\, \U1/N_2151\, \U1/N_2152\, \U1/N_698\, 
        \U1/N_2153\, \U1/N_2154\, \U1/N_700\, \U1/N_2155\, 
        \U1/N_2156\, \U1/N_702\, \U1/N_704\, \U1/N_2159\, 
        \U1/N_2160\, \U1/N_706\, \U1/N_708\, \U1/N_2163\, 
        \U1/N_2164\, \U1/N_333\, \U1/N_329\, \U1/N_327\, 
        \U1/N_325\, \U1/N_323\, \U1/N_321\, \U1/N_319\, 
        \U1/N_317\, \U1/N_1816\, \U1/N_1815\, \U1/N_1814\, 
        \U1/N_724\, \U1/N_296\, \U1/N_284\, \U1/N_2197\, 
        \U1/N_2198\, \U1/N_278\, \U1/N_2199\, \U1/N_2200\, 
        \U1/N_272\, \U1/N_266\, \U1/N_1812\, \U1/N_2205\, 
        \U1/N_2206\, \U1/N_1811\, \U1/N_1810\, \U1/N_1808\, 
        \U1/N_1807\, \U1/N_154\, \U1/N_2217\, \U1/N_2218\, 
        \U1/N_1806\, \U1/N_1805\, \U1/N_742\, \U1/N_1801\, 
        \U1/N_1800\, \U1/N_1799\, \U1/N_2231\, \U1/N_2232\, 
        \U1/N_1798\, \U1/N_130\, \U1/N_751\, \U1/N_1797\, 
        \U1/N_124\, \U1/N_122\, \U1/N_1796\, \U1/N_1795\, 
        \U1/N_2247\, \U1/N_2248\, \U1/N_1794\, \U1/N_763\, 
        \U1/N_1792\, \U1/N_2255\, \U1/N_2256\, \U1/N_1791\, 
        \U1/N_1790\, \U1/N_1789\, \U1/N_1788\, \U1/N_772\, 
        \U1/N_1787\, \U1/N_1786\, \U1/N_2269\, \U1/N_2270\, 
        \U1/N_1785\, \U1/N_1784\, \U1/N_1783\, \U1/N_2275\, 
        \U1/N_2276\, \U1/N_1782\, \U1/N_1779\, \U1/N_1610\, 
        \U1/N_1778\, \U1/N_1777\, \U1/N_1776\, \U1/N_1775\, 
        \U1/N_2291\, \U1/N_2292\, \U1/N_787\, \U1/N_789\, 
        \U1/N_2295\, \U1/N_2296\, \U1/pr_state_RNO[3]_net_1\, 
        \U1/N_858\, \U1/N_158\, \U1/N_17\, \U1/N_91\, \U1/N_70\, 
        \U1/N_51\, \U1/N271\, \U1/N270\, \U1/N315\, \U1/N313\, 
        \U1/cnt_daly_n9\, \U1/cnt_daly_n10\, \U1/cnt_n2_net_1\, 
        \U1/cnt_63_0_net_1\, \U1/data_filter_4[12]\, 
        \U1/data_filter_4[13]\, \U1/N200\, \U1/N201\, \U1/N203\, 
        \U1/N204\, \U1/N197\, \U1/N240\, \U1/N241\, \U1/N267\, 
        \U1/N244\, \U1/N248\, \U1/I71_un1_Y\, \U1/N188\, 
        \U1/N247\, \U1/N186\, \U1/N183\, \U1/N195\, \U1/N179\, 
        \U1/N182\, \U1/N180\, \U1/N185\, \U1/N191\, \U1/N194\, 
        \U1/data_all_3[175]\, \U1/data_all_3[174]\, 
        \U1/data_all_3[79]\, \U1/data_all_3[78]\, 
        \U1/data_all_3[47]\, \U1/data_all_3[46]\, 
        \U1/data_all_3[159]\, \U1/data_all_3[158]\, 
        \U1/data_all_3[31]\, \U1/data_all_3[30]\, 
        \U1/data_all_3[95]\, \U1/data_all_3[94]\, 
        \U1/data_all_3[15]\, \U1/data_all_3[14]\, \U1/N_18\, 
        \U1/N_1781\, \U1/N_867\, \U1/N_834\, \U1/N_1093\, 
        \U1/N_1094\, \U1/N_1092\, \U1/N_793\, \U1/N_1838\, 
        \U1/N_872\, \U1/N_1415\, \U1/cnt_n1_net_1\, \U1/N_859\, 
        \U1/cnt_daly_n12\, \U1/cnt_daly_n11\, \U1/N_42\, 
        \U1/N_1090\, \U1/delay_channel1_net_1\, 
        \U1/pr_state_ns[3]\, \U1/N207\, \U1/N_260\, \U1/N_263\, 
        \U1/cnt_receive_over_1_sqmuxa_net_1\, \U1/N_3\, 
        \U0/conver_ris2_i\, \U0/conver_ris2_net_1\, 
        \U0/pr_state_ns_a4_2[1]\, \U0/pr_state[0]_net_1\, 
        \U0/cnt_rc[3]_net_1\, \U0/cnt_rc[1]_net_1\, 
        \U0/cnt_rc[2]_net_1\, \U0/cnt_rc[0]_net_1\, 
        \U0/cnt_rc_7_0_net_1\, \U0/pr_state[4]_net_1\, 
        \U0/pr_state_ns[1]\, \U0/cnt_rc_n2_net_1\, \U0/N_130\, 
        \U0/data_ad_4[0]\, \U0/pr_state[5]_net_1\, 
        \U0/data_ad_4[1]\, \U0/data_ad_4[2]\, \U0/data_ad_4[3]\, 
        \U0/data_ad_4[4]\, \U0/data_ad_4[5]\, \U0/data_ad_4[6]\, 
        \U0/data_ad_4[7]\, \U0/data_ad_4[9]\, \U0/data_ad_4[11]\, 
        \U0/N_138\, \U0/pr_state[2]_net_1\, \U0/un1_pr_state_5\, 
        \U0/N_137\, \U0/pr_state[1]_net_1\, \U0/cnt_rc_n3_net_1\, 
        \U0/N_59\, \U0/cnt_rc_n1_net_1\, \U0/N_164\, 
        \U0/pr_state_RNO_0[0]_net_1\, \U0/N_143\, 
        \U0/pr_state_RNO[2]_net_1\, \U0/pr_state[3]_net_1\, 
        \U0/sts_ris_i_0\, \U0/pr_state_ns[2]\, 
        \U0/pr_state_ns[0]\, \U0/conver_ris_i_0\, \U0/N_144\, 
        \U0/N_136\, \U0/N_135\, \U0/data_ad_4[10]\, 
        \U0/data_ad_4[8]\, \U0/conver_ris_1\, 
        \U0/conver_ris3_i_0\, \U0/sts_ris_2\, \U0/sts_ris3_net_1\, 
        \U0/sts_ris2_net_1\, \U0/sts_ris1_net_1\, 
        \U0/conver_ris1_net_1\, \U5/cnt_0[2]_net_1\, \U5/cnt_n2\, 
        \U5/pr_state[0]_net_1\, \U5/cnt[1]_net_1\, \U5/cnt_0[1]\, 
        \U5/cnt[0]_net_1\, \U5/cnt_0[0]\, 
        \U5/pr_state_ns_0_i_0[0]\, \U5/pr_state_ns_0_i_a4_0_0[0]\, 
        \U5/N_7\, \U5/m7_1\, \U5/cnt[3]_net_1\, \U5/cnt[4]_net_1\, 
        \U5/cnt[2]_net_1\, \U5/pr_state[1]_net_1\, \U5/N_6\, 
        \U5/N_138_mux\, \U5/pr_state_RNO[1]_net_1\, \U5/N_339\, 
        \U5/N_340\, \U5/N_341\, \U5/N_343\, \U5/N_344\, 
        \U5/N_345\, \U5/N_346\, \U5/N_347\, \U5/N_348\, 
        \U5/N_349\, \U5/N_351\, \U5/N_352\, \U5/N_353\, 
        \U5/N_354\, \U5/N_355\, \U5/N_356\, \U5/N_357\, 
        \U5/N_359\, \U5/N_360\, \U5/N_361\, \U5/N_362\, 
        \U5/N_363\, \U5/N_364\, \U5/N_365\, \U5/N_367\, 
        \U5/N_368\, \U5/N_369\, \U5/N_370\, \U5/N_371\, 
        \U5/N_372\, \U5/N_373\, \U5/N_374\, \U5/N_375\, 
        \U5/N_377\, \U5/N_378\, \U5/N_379\, \U5/N_380\, 
        \U5/N_381\, \U5/N_382\, \U5/N_383\, \U5/N_385\, 
        \U5/N_386\, \U5/N_387\, \U5/N_388\, \U5/N_389\, 
        \U5/N_390\, \U5/N_391\, \U5/N_393\, \U5/N_394\, 
        \U5/N_395\, \U5/N_396\, \U5/N_397\, \U5/N_398\, 
        \U5/N_399\, \U5/N_401\, \U5/N_402\, \U5/N_403\, 
        \U5/N_404\, \U5/N_405\, \U5/N_406\, \U5/N_407\, 
        \U5/N_409\, \U5/N_410\, \U5/N_411\, \U5/N_413\, 
        \U5/N_414\, \U5/N_415\, \U5/N_417\, \U5/N_418\, 
        \U5/N_419\, \U5/N_421\, \U5/N_422\, \U5/N_423\, 
        \U5/N_425\, \U5/N_426\, \U5/N_427\, \U5/N_429\, 
        \U5/N_430\, \U5/N_433\, \U5/N_434\, \U5/N_435\, 
        \U5/N_436\, \U5/N_437\, \U5/N_438\, \U5/N_441\, 
        \U5/N_442\, \U5/N_443\, \U5/N_444\, \U5/N_445\, 
        \U5/N_446\, \U5/N_449\, \U5/N_450\, \U5/N_451\, 
        \U5/N_452\, \U5/N_453\, \U5/N_454\, \U5/N_457\, 
        \U5/N_458\, \U5/N_459\, \U5/N_460\, \U5/N_461\, 
        \U5/N_463\, \U5/N_464\, \U5/N_465\, \U5/N_466\, 
        \U5/N_467\, \U5/N_468\, \U5/N_469\, \U5/N_471\, 
        \U5/N_472\, \U5/N_473\, \U5/N_474\, \U5/N_475\, 
        \U5/N_476\, \U5/N_477\, \U5/N_478\, \U5/N_479\, 
        \U5/N_481\, \U5/N_482\, \U5/N_483\, \U5/N_484\, 
        \U5/N_485\, \U5/N_486\, \U5/N_487\, \U5/N_488\, 
        \U5/N_392\, \U5/N_400\, \U5/N_489\, \U5/N_490\, 
        \U5/N_491\, \U5/N_493\, \U5/N_494\, \U5/N_495\, 
        \U5/N_497\, \U5/N_498\, \U5/N_499\, \U5/N_501\, 
        \U5/N_502\, \U5/N_503\, \U5/N_431\, \U5/N_505\, 
        \U5/N_506\, \U5/N_507\, \U5/N_508\, \U5/N_509\, 
        \U5/N_510\, \U5/N_513\, \U5/N_514\, \U5/N_515\, 
        \U5/N_516\, \U5/N_517\, \U5/N_519\, \U5/N_520\, 
        \U5/N_521\, \U5/N_522\, \U5/N_523\, \U5/N_525\, 
        \U5/N_526\, \U5/N_527\, \U5/N_529\, \U5/N_25_0\, 
        \U5/N_26_0\, \U5/N_27_0\, \U5/N_530\, 
        \U5/un58_data_send[7]\, \U5/i58_mux\, \U5/N_32_0\, 
        \U5/N_33_0\, \U5/N_34_0\, \U5/N_531\, 
        \U5/un58_data_send[6]\, \U5/i71_mux\, \U5/N_46_0\, 
        \U5/N_455\, \U5/N_47_0\, \U5/N_511\, \U5/N_48_0\, 
        \U5/N_533\, \U5/un58_data_send[4]\, \U5/i67_mux\, 
        \U5/N_53_0\, \U5/N_54_0\, \U5/N_55_0\, \U5/N_534\, 
        \U5/un58_data_send[3]\, \U5/i65_mux\, \U5/N_60_0\, 
        \U5/N_61_0\, \U5/N_62_0\, \U5/N_535\, 
        \U5/un58_data_send[2]\, \U5/i63_mux\, \U5/N_67_0\, 
        \U5/N_68\, \U5/N_74\, \U5/N_75\, \U5/N_76\, \U5/N_537\, 
        \U5/un58_data_send[0]\, \U5/i59_mux\, \U5/N_538\, 
        \U5/N_518\, \U5/N_78\, \U5/un1_pr_state_1\, \U5/N_39_0\, 
        \U5/N_456\, \U5/N_432\, \U5/N_424\, \U5/N_416\, 
        \U5/N_408\, \U5/N_376\, \U5/N_384\, \U5/N_440\, 
        \U5/N_448\, \U5/N_480\, \U5/N_496\, \U5/N_504\, 
        \U5/N_512\, \U5/N_528\, \U5/N_40_0\, \U5/N_41_0\, 
        \U5/N_116\, \U5/un58_data_send[5]\, \U5/i69_mux\, 
        \U5/i61_mux\, \U5/N_524\, \U5/N_536\, \U5/N_492\, 
        \U5/N_500\, \U5/un58_data_send[1]\, \U5/N_69\, 
        \U5/N_21_0\, \U5/cnt_n1\, \U5/N_10_0\, \U5/cnt_n3\, 
        \U5/N_11_0\, \U5/cnt_n4\, \U5/N_12_0\, \U5/N_462\, 
        \U5/N_470\, \U5/N_439\, \U5/N_447\, \U5/N_420\, 
        \U5/N_428\, \U5/N_412\, \U5/N_358\, \U5/N_366\, 
        \U5/N_342\, \U5/N_350\, \data_in_pad[8]/U0/NET1\, 
        \data_in_pad[10]/U0/NET1\, \ce_pad/U0/NET1\, 
        \ce_pad/U0/NET2\, \addr_pad[0]/U0/NET1\, 
        \addr_pad[0]/U0/NET2\, \rc_pad/U0/NET1\, \rc_pad/U0/NET2\, 
        \data_in_pad[6]/U0/NET1\, \data_in_pad[7]/U0/NET1\, 
        \data_in_pad[5]/U0/NET1\, \data_in_pad[11]/U0/NET1\, 
        \sys_clk_pad/U0/NET1\, \sys_rest_pad/U0/NET1\, 
        \data_in_pad[3]/U0/NET1\, \data_in_pad[4]/U0/NET1\, 
        \addr_pad[3]/U0/NET1\, \addr_pad[3]/U0/NET2\, 
        \data_in_pad[9]/U0/NET1\, \sts_pad/U0/NET1\, 
        \rx_uart_pad/U0/NET1\, \data_in_pad[1]/U0/NET1\, 
        \addr_pad[2]/U0/NET1\, \addr_pad[2]/U0/NET2\, 
        \data_in_pad[0]/U0/NET1\, \tx_uart_pad/U0/NET1\, 
        \tx_uart_pad/U0/NET2\, \cs_pad/U0/NET1\, \cs_pad/U0/NET2\, 
        \data_in_pad[2]/U0/NET1\, \addr_pad[1]/U0/NET1\, 
        \addr_pad[1]/U0/NET2\, \VCC\, AFLSDF_VCC, AFLSDF_GND
         : std_logic;
    signal GND_power_net1 : std_logic;
    signal VCC_power_net1 : std_logic;

begin 

    AFLSDF_GND <= GND_power_net1;
    \GND\ <= GND_power_net1;
    \VCC\ <= VCC_power_net1;
    AFLSDF_VCC <= VCC_power_net1;

    \U1/data_all_RNO_0[37]\ : AO1C
      port map(A => \data_all[37]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m283_i_0_0\);
    
    \U1/data_all_3_0_0_i_o2_0_0[92]\ : OR2
      port map(A => \U1/N_826\, B => \U1/N_821\, Y => 
        \U1/N_834_0\);
    
    \U2/cnt_RNILL7J[4]\ : NOR3B
      port map(A => \U2/cnt[5]_net_1\, B => \U2/un1_cnt_1\, C => 
        \U2/cnt[4]_net_1\, Y => \U2/tx_uart36_7\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I46_Y\ : AO1
      port map(A => \U1/N242\, B => \U1/N239\, C => \U1/N238\, Y
         => \U1/N265\);
    
    \U5/data_send_RNO_23[2]\ : MX2
      port map(A => \data_all[146]\, B => \data_all[154]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_413\);
    
    \U2/parity_check_RNO_9\ : XA1A
      port map(A => \U2/parity_check_net_1\, B => \data_send[4]\, 
        C => \U2/parity_check_5_sqmuxa\, Y => \U2/N_121\);
    
    \U1/m146_i_0_o2\ : OR2
      port map(A => \U1/m146_i_0_o2_1\, B => \U1/N_817\, Y => 
        \U1/N_838\);
    
    \U1/data_all_RNO_1[219]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_840\, 
        Y => \U1/N_1018\);
    
    \U1/data_all[6]\ : DFN1E0C0
      port map(D => \U1/N_250\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[6]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I79_Y\ : OR3
      port map(A => \U1/I79_un1_Y\, B => 
        \U1/ADD_14x14_fast_I79_Y_0\, C => \U1/I64_un1_Y\, Y => 
        \U1/N319\);
    
    \U5/data_send_RNO_8[3]\ : MX2
      port map(A => \U5/N_374\, B => \U5/N_382\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_478\);
    
    \U1/data_all_RNO[183]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[183]\, Y => \U1/N_407\);
    
    \U1/data_all[28]\ : DFN1E0C0
      port map(D => \U1/N_765\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[28]\);
    
    \U0/data_ad_RNO[2]\ : NOR2A
      port map(A => \data_in_c[2]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[2]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I37_Y\ : NOR2B
      port map(A => \U1/N229\, B => \U1/N233\, Y => \U1/N256\);
    
    \U1/data_all_RNO[86]\ : OA1B
      port map(A => \U1/N_834_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[86]\, Y => \U1/N_205\);
    
    \U1/data_all_RNO[180]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[180]\, Y => \U1/N_401\);
    
    \U5/data_send_RNO_18[5]\ : MX2
      port map(A => \data_all[69]\, B => \data_all[77]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_376\);
    
    \data_in_pad[8]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[8]/U0/NET1\, Y => 
        \data_in_c[8]\);
    
    \U3/data_recive_RNO_2[3]\ : NOR3A
      port map(A => \U3/m36_1\, B => \U3/cnt[0]_net_1\, C => 
        \U3/cnt[1]_net_1\, Y => \U3/m36_4\);
    
    \U1/data_all_RNO_1[202]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_839\, 
        Y => \U1/N_926\);
    
    \U2/cnt_c7\ : NOR2B
      port map(A => \U2/cnt_c6_net_1\, B => \U2/cnt[7]_net_1\, Y
         => \U2/cnt_c7_net_1\);
    
    \U1/data_all[125]\ : DFN1E0C0
      port map(D => \U1/N_390\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[125]\);
    
    \U5/pr_state_RNO_0[0]\ : MX2
      port map(A => \U5/pr_state_ns_0_i_a4_0_0[0]\, B => \U5/N_7\, 
        S => \U5/pr_state[0]_net_1\, Y => 
        \U5/pr_state_ns_0_i_0[0]\);
    
    \U2/cnt_RNI3KRS[1]\ : NOR3C
      port map(A => \U2/un1_cnt_3\, B => \U2/N_165\, C => 
        \U2/N_163\, Y => \U2/tx_uart33_0_a2_0_2\);
    
    \U1/data_all[148]\ : DFN1E0C0
      port map(D => \U1/N_124\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[148]\);
    
    \U5/data_send_RNO_4[1]\ : MX2C
      port map(A => \U5/N_492\, B => \U5/N_500\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_536\);
    
    \U1/data_all_RNO[165]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m179_i_0_0\, Y => \U1/N_317\);
    
    \U1/data_all[168]\ : DFN1E0C0
      port map(D => \U1/N_323\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[168]\);
    
    \U2/parity_check\ : DFN1E0P0
      port map(D => \U2/parity_check_10_iv\, CLK => sys_clk_c, 
        PRE => sys_rest_c, E => \U2/parity_check_0_sqmuxa\, Q => 
        \U2/parity_check_net_1\);
    
    \U1/data_all_RNO[42]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2199\, C
         => \U1/N_2200\, Y => \U1/N_278\);
    
    \U1/data_all_RNO_0[97]\ : AO1C
      port map(A => \data_all[97]\, B => \U1/N_829_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[97]\);
    
    \U1/data_all_RNO_0[8]\ : AO1C
      port map(A => \data_all[8]\, B => \U1/N_835\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[8]\);
    
    \U1/data_all_RNO_0[103]\ : AO1C
      port map(A => \data_all[103]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[103]\);
    
    \U3/data_recive_RNO_3[7]\ : NOR2A
      port map(A => \U3/cnt[8]_net_1\, B => \U3/cnt[1]_net_1\, Y
         => \U3/m22_1\);
    
    \U3/data_recive_RNO_3[4]\ : NOR2A
      port map(A => \U3/cnt[3]_net_1\, B => \U3/cnt[1]_net_1\, Y
         => \U3/m53_2\);
    
    \U1/data_all[157]\ : DFN1E0C0
      port map(D => \U1/N_742\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[157]\);
    
    \U3/data_recive[0]\ : DFN1C0
      port map(D => \U3/data_recive_12[0]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[0]\);
    
    \U1/data_all_RNO_0[107]\ : AO1C
      port map(A => \data_all[107]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[107]\);
    
    \U5/data_send_RNO_26[7]\ : MX2
      port map(A => \data_all[199]\, B => \data_all[207]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_442\);
    
    \U1/data_all_RNO_0[35]\ : AO1C
      port map(A => \data_all[35]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m289_i_0_0\);
    
    \U1/cnt_daly_RNI1GVQ[6]\ : NOR2A
      port map(A => \U1/cnt_daly[7]_net_1\, B => 
        \U1/cnt_daly[6]_net_1\, Y => \U1/m61_0_i_a3_1_5\);
    
    \U0/cnt_rc_7_0\ : NOR2A
      port map(A => \U0/cnt_rc[2]_net_1\, B => 
        \U0/pr_state[4]_net_1\, Y => \U0/cnt_rc_7_0_net_1\);
    
    \U5/data_send_RNO_12[1]\ : MX2
      port map(A => \U5/N_436\, B => \U5/N_444\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_508\);
    
    \U1/data_all_RNO[215]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1021\, C
         => \U1/N_1022\, Y => \U1/N_178\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I9_P0N\ : OR2
      port map(A => \data_ad[9]\, B => \U1/data_filter[9]_net_1\, 
        Y => \U1/N204\);
    
    \U2/cnt[4]\ : DFN1C0
      port map(D => \U2/cnt_n4_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[4]_net_1\);
    
    \U1/data_all[22]\ : DFN1E0C0
      port map(D => \U1/N_772\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[22]\);
    
    \U5/data_send_RNO_13[6]\ : NOR2A
      port map(A => \U5/N_457\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_32_0\);
    
    \U1/data_all_RNO_0[86]\ : AO1C
      port map(A => \data_all[86]\, B => \U1/N_834_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[86]\);
    
    \U1/data_all_RNO[118]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[118]\, Y => \U1/N_376\);
    
    \U1/cnt_receive_over\ : DFN1E0C0
      port map(D => addr_over_i, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/cnt_receive_over_1_sqmuxa_net_1\, Q
         => \U1/cnt_receive_over_net_1\);
    
    \U1/data_all_RNO[66]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/m246_i_0_0\, Y => \U1/N_167\);
    
    \U0/data_ad[9]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[9]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[9]\);
    
    \U1/data_all_RNO_0[89]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[89]\, Y => 
        \U1/N_2133\);
    
    \U1/data_all_3_0_a2_i_0_o2[239]\ : OR2
      port map(A => \U1/m146_i_0_o2_1\, B => \U1/N_818\, Y => 
        \U1/N_837\);
    
    \U1/cnt_daly[12]\ : DFN1E0C0
      port map(D => \U1/cnt_daly_n12\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => 
        \U1/cnt_daly[12]_net_1\);
    
    \U5/pr_state_RNO_1[0]\ : OA1C
      port map(A => vld_whole, B => send_whole_over, C => 
        \U5/pr_state[1]_net_1\, Y => 
        \U5/pr_state_ns_0_i_a4_0_0[0]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I33_Y\ : NOR2B
      port map(A => \U1/N180\, B => \U1/N183\, Y => \U1/N249\);
    
    \U1/m103_i_o2_0_o2\ : OR2
      port map(A => \U1/m103_i_o2_0_o2_0_net_1\, B => \U1/N_818\, 
        Y => \U1/N_839\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I78_Y_0\ : AO1
      port map(A => \U1/N236\, B => \U1/N233\, C => \U1/N232\, Y
         => \U1/ADD_14x14_fast_I78_Y_0\);
    
    \U1/data_all_RNO[175]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_838\, C
         => \data_all[175]\, Y => \U1/data_all_3[175]\);
    
    \U5/data_send_RNO_15[4]\ : MX2
      port map(A => \data_all[20]\, B => \data_all[28]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_351\);
    
    \U5/data_send_RNO_14[5]\ : MX2
      port map(A => \data_all[5]\, B => \data_all[13]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_344\);
    
    \U1/data_all_RNO[52]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[52]\, Y => \U1/N_694\);
    
    \U2/cnt_RNI1J3G1[1]\ : NOR2B
      port map(A => \U2/tx_uart33_0_a2_0_2\, B => \U2/N_171\, Y
         => \U2/N_197\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I50_Y\ : AO1
      port map(A => \U1/N246\, B => \U1/N243\, C => \U1/N242\, Y
         => \U1/N269\);
    
    \U5/data_send_RNO_12[4]\ : MX2
      port map(A => \U5/N_439\, B => \U5/N_447\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_511\);
    
    \U1/data_all_RNO[136]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/m199_0_i_0\, Y => \U1/N_103\);
    
    \U5/data_send_RNO_11[5]\ : MX2
      port map(A => \U5/N_424\, B => \U5/N_432\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_504\);
    
    \U2/cnt_RNIUI2J1[10]\ : NOR2B
      port map(A => \U2/N_153\, B => \U2/N_127\, Y => \U2/N_173\);
    
    \U3/cnt_4[5]\ : XA1
      port map(A => \U3/N_8\, B => \U3/cnt[5]_net_1\, C => 
        \U3/recive_net_1\, Y => \U3/cnt_4[5]_net_1\);
    
    \U1/data_all_RNO[155]\ : OA1B
      port map(A => \U1/N_842\, B => \U1/data_filter[11]_net_1\, 
        C => \U1/m83_1_i_0_0\, Y => \U1/N_1801\);
    
    \U0/conver_ris1\ : DFN1C0
      port map(D => conver_top, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U0/conver_ris1_net_1\);
    
    \U2/parity_check_RNO_8\ : XA1A
      port map(A => \U2/parity_check_net_1\, B => \data_send[0]\, 
        C => \U2/parity_check_1_sqmuxa\, Y => \U2/N_116\);
    
    \U1/data_all_RNO_0[13]\ : AO1C
      port map(A => \data_all[13]\, B => \U1/N_835_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[13]\);
    
    \U4/pr_state_RNIR2CG[0]\ : NOR2A
      port map(A => \U4/pr_state[0]_net_1\, B => \addr_c[0]\, Y
         => \U4/N_20\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I89_Y\ : XOR3
      port map(A => \U1/data_filter[1]_net_1\, B => \data_ad[1]\, 
        C => \U1/N176\, Y => \U1/un2_data_filter[1]\);
    
    \U1/data_all_RNO_0[145]\ : NOR2A
      port map(A => \U1/N_842\, B => \data_all[145]\, Y => 
        \U1/N_2247\);
    
    \U1/data_all[170]\ : DFN1E0C0
      port map(D => \U1/N_327\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[170]\);
    
    \U5/data_send_RNO_18[7]\ : MX2
      port map(A => \data_all[71]\, B => \data_all[79]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_378\);
    
    \U1/data_all_RNO_0[1]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[1]\, Y => 
        \U1/N_1098\);
    
    \U1/data_all[3]\ : DFN1E0C0
      port map(D => \U1/N_258\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[3]\);
    
    \U1/data_all_RNO[196]\ : OA1B
      port map(A => \U1/N_839\, B => \U1/data_filter[4]_net_1\, C
         => \U1/m133_i_0_0\, Y => \U1/N_203\);
    
    \U1/data_all_RNO[148]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/m106_0_i_0_0\, Y => \U1/N_124\);
    
    \U1/data_all[181]\ : DFN1E0C0
      port map(D => \U1/N_403\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[181]\);
    
    \U5/data_send_RNO_5[6]\ : MX2
      port map(A => \U5/N_513\, B => \U5/N_32_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_33_0\);
    
    \U1/data_all[21]\ : DFN1E0C0
      port map(D => \U1/N_1787\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[21]\);
    
    \U4/addr_RNIK2EN[3]\ : NOR3
      port map(A => \addr_c[2]\, B => \addr_c[3]\, C => 
        \addr_c[1]\, Y => \U4.N_31\);
    
    \U1/data_all[27]\ : DFN1E0C0
      port map(D => \U1/N_1792\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[27]\);
    
    \U5/data_send_RNO_21[2]\ : MX2
      port map(A => \data_all[114]\, B => \data_all[122]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_397\);
    
    \U3/data_recive[6]\ : DFN1C0
      port map(D => \U3/data_recive_12[6]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[6]\);
    
    \U2/cnt_RNIH1K9_2[8]\ : NOR2
      port map(A => \U2/cnt[8]_net_1\, B => \U2/cnt[5]_net_1\, Y
         => \U2/N_166\);
    
    \U1/data_all_RNO_0[72]\ : AO1C
      port map(A => \data_all[72]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m228_i_0_0\);
    
    \U1/m206_i_0_o2\ : OR2
      port map(A => \U1/N_826\, B => \U1/N_819\, Y => \U1/N_833\);
    
    \U1/data_all_RNO_1[91]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_834\, 
        Y => \U1/N_2132\);
    
    \U1/data_all_RNO_0[235]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[235]\, Y => 
        \U1/N_909\);
    
    \U1/data_all_RNO[167]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/m173_i_0_0\, Y => \U1/N_321\);
    
    \U1/data_all_RNO_0[45]\ : AO1C
      port map(A => \data_all[45]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m258_i_0_0\);
    
    \U1/data_all[132]\ : DFN1E0C0
      port map(D => \U1/N_245\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[132]\);
    
    \U1/data_all_RNO[232]\ : OA1B
      port map(A => \U1/N_837_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/m82_0_i_0_0\, Y => \U1/N_221\);
    
    \U2/cnt_RNI7DUF2_1[10]\ : NOR2B
      port map(A => \U2/N_192\, B => \U2/N_168\, Y => 
        \U2/parity_check_8_sqmuxa\);
    
    \U2/parity_check_RNO_5\ : XOR2
      port map(A => \data_send[2]\, B => \U2/parity_check_net_1\, 
        Y => \U2/N_68_i\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I99_Y_0\ : XOR2
      port map(A => \data_ad[11]\, B => 
        \U1/data_filter[11]_net_1\, Y => 
        \U1/ADD_14x14_fast_I99_Y_0\);
    
    \U2/tx_uart_RNO_1\ : AO1
      port map(A => \U2/parity_check_6_sqmuxa\, B => 
        \data_send[5]\, C => \U2/tx_uart_11_iv_2\, Y => 
        \U2/tx_uart_11_iv_6\);
    
    \U5/cnt_RNO_0[4]\ : NOR2B
      port map(A => \U5/N_11_0\, B => \U5/cnt[3]_net_1\, Y => 
        \U5/N_12_0\);
    
    \U2/cnt_RNIETQ61[0]\ : NOR2B
      port map(A => \U2/N_165\, B => \U2/N_154\, Y => 
        \U2/tx_uart27_0_a2_3\);
    
    \U5/data_send_RNO_5[5]\ : MX2
      port map(A => \U5/N_512\, B => \U5/N_39_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_40_0\);
    
    \U5/data_send_RNO_18[3]\ : MX2
      port map(A => \data_all[67]\, B => \data_all[75]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_374\);
    
    \U1/data_all_RNO[133]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[133]\, Y => \U1/N_1836\);
    
    \U1/data_all_RNO_0[179]\ : AO1C
      port map(A => \data_all[179]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[179]\);
    
    \U3/cnt_RNIS0VF[10]\ : NOR2B
      port map(A => \U3/cnt[10]_net_1\, B => \U3/cnt[5]_net_1\, Y
         => \U3/m22_0\);
    
    \U5/pr_state[0]\ : DFN1C0
      port map(D => \U5/N_6\, CLK => sys_clk_c, CLR => sys_rest_c, 
        Q => \U5/pr_state[0]_net_1\);
    
    \U1/data_all_RNO_0[176]\ : AO1C
      port map(A => \data_all[176]\, B => \U1/N_844_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[176]\);
    
    \U1/data_all_RNO[130]\ : OA1B
      port map(A => \U1/N_841\, B => \U1/data_filter[2]_net_1\, C
         => \U1/m205_0_i_0\, Y => \U1/N_107\);
    
    \U1/data_all[144]\ : DFN1E0C0
      port map(D => \U1/N_1794\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[144]\);
    
    \U3/cnt_RNIICDP[4]\ : NOR3B
      port map(A => \U3/cnt[4]_net_1\, B => \U3/cnt[3]_net_1\, C
         => \U3/cnt[2]_net_1\, Y => \U3/m11_6\);
    
    \U1/pr_state_RNIPCN11[4]\ : NOR3
      port map(A => \U1/pr_state_0[7]_net_1\, B => 
        \U1/pr_state[4]_net_1\, C => \U1/pr_state[5]_net_1\, Y
         => \U1/N_1094\);
    
    \U3/data_recive_RNO_3[5]\ : NOR2A
      port map(A => \U3/cnt[1]_net_1\, B => \U3/cnt[3]_net_1\, Y
         => \U3/m47_2\);
    
    \U1/data_all_RNO_0[172]\ : AO1C
      port map(A => \data_all[172]\, B => \U1/N_838_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m156_i_0_0\);
    
    \U1/data_all_RNO[45]\ : OA1B
      port map(A => \U1/N_832\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m258_i_0_0\, Y => \U1/N_296\);
    
    \U1/data_all[191]\ : DFN1E0C0
      port map(D => \U1/N_51\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[191]\);
    
    \U1/data_all[164]\ : DFN1E0C0
      port map(D => \U1/N_315\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[164]\);
    
    \U1/data_all_RNO_0[149]\ : AO1C
      port map(A => \data_all[149]\, B => \U1/N_842\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m103_0_i_0_0\);
    
    \U5/data_send_RNO_0[0]\ : MX2C
      port map(A => \U5/N_515\, B => \U5/N_523\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i59_mux\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I76_un1_Y_0\ : NOR2B
      port map(A => \U1/N256\, B => \U1/N264\, Y => 
        \U1/ADD_14x14_fast_I76_un1_Y_0\);
    
    \U1/data_all_RNO_1[2]\ : NOR2
      port map(A => \U1/data_filter[2]_net_1\, B => \U1/N_835\, Y
         => \U1/N_982\);
    
    \U1/data_all_RNO_0[146]\ : AO1C
      port map(A => \data_all[146]\, B => \U1/N_842\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m112_1_i_0_0\);
    
    \U1/data_all_RNO_0[178]\ : AO1C
      port map(A => \data_all[178]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[178]\);
    
    \U1/data_all_RNO[193]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[1]_net_1\, 
        C => \U1/m142_0_i_0\, Y => \U1/N_96\);
    
    \U1/data_all_RNO[177]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[1]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[177]\, Y => \U1/N_395\);
    
    \U5/data_send_RNO_17[0]\ : MX2
      port map(A => \data_all[48]\, B => \data_all[56]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_363\);
    
    \U1/data_filter_RNO[5]\ : OA1C
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/un2_data_filter[5]\, C => \U1/m54_0_0_0\, Y => 
        \U1/N_55_0\);
    
    \U5/cnt_RNO[1]\ : XA1
      port map(A => \U5/cnt[0]_net_1\, B => \U5/cnt[1]_net_1\, C
         => \U5/pr_state[1]_net_1\, Y => \U5/cnt_n1\);
    
    \U1/data_all_RNO_1[89]\ : NOR2
      port map(A => \U1/data_filter[9]_net_1\, B => \U1/N_834\, Y
         => \U1/N_2134\);
    
    \U1/data_all_RNO[190]\ : NOR3C
      port map(A => \data_all[190]\, B => \U1/pr_state[2]_net_1\, 
        C => \U1/N_844\, Y => \U1/N_53\);
    
    \U2/cnt_RNICSJ9_0[2]\ : NOR2A
      port map(A => \U2/cnt[6]_net_1\, B => \U2/cnt[2]_net_1\, Y
         => \U2/tx_uart37_3\);
    
    \U2/cnt[3]\ : DFN1C0
      port map(D => \U2/cnt_n3_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[3]_net_1\);
    
    \U1/data_all_RNO[23]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/m144_0_i_0_0\, Y => \U1/N_1788\);
    
    \U1/data_all_RNO[224]\ : OA1B
      port map(A => \U1/N_837_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[224]\, Y => \U1/N_34\);
    
    \U5/data_send_RNO_26[4]\ : MX2
      port map(A => \data_all[196]\, B => \data_all[204]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_439\);
    
    \U3/data_recive_RNO_1[1]\ : NOR3C
      port map(A => \U3/m27_2\, B => \U3/m27_1\, C => 
        \U3/N_125_mux\, Y => \U3/data_recive24\);
    
    \U1/data_all[117]\ : DFN1E0C0
      port map(D => \U1/N_374\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[117]\);
    
    \U1/data_filter_RNO[13]\ : XA1
      port map(A => \U1/data_filter[13]_net_1\, B => \U1/N313\, C
         => \U1/pr_state_0[5]_net_1\, Y => \U1/data_filter_4[13]\);
    
    \U1/data_all_RNO_0[148]\ : AO1C
      port map(A => \data_all[148]\, B => \U1/N_842_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m106_0_i_0_0\);
    
    \U1/data_all[122]\ : DFN1E0C0
      port map(D => \U1/N_384\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[122]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I3_G0N\ : NOR2B
      port map(A => \data_ad[3]\, B => \U1/data_filter[3]_net_1\, 
        Y => \U1/N185\);
    
    \U1/data_all_RNO[157]\ : OA1B
      port map(A => \U1/N_842\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m79_0_i_i_0\, Y => \U1/N_742\);
    
    \U1/data_all_3_0_a2_i_0_o2_2[239]\ : OR2A
      port map(A => \U1/I_7_0\, B => \U1/OVER\, Y => \U1/N_818\);
    
    \U1/data_all_RNO[38]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/m280_i_0_0\, Y => \U1/N_1811\);
    
    \U1/data_all_RNO[217]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1019\, C
         => \U1/N_1020\, Y => \U1/N_174\);
    
    \U1/data_all[74]\ : DFN1E0C0
      port map(D => \U1/N_183\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[74]\);
    
    \U1/m79_0_i_i_o2_0\ : OR3A
      port map(A => \U1/I_9_0\, B => \addr_c_0[0]\, C => 
        \U1/I_5_0\, Y => \U1/m79_0_i_i_o2_0_net_1\);
    
    \U1/m79_0_i_i_o2\ : OR2
      port map(A => \U1/m79_0_i_i_o2_0_net_1\, B => \U1/N_817\, Y
         => \U1/N_842\);
    
    \U1/data_filter[8]\ : DFN1E0C0
      port map(D => \U1/N_39\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[8]_net_1\);
    
    \data_in_pad[0]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[0]/U0/NET1\, Y => 
        \data_in_c[0]\);
    
    \U2/cnt_RNI6VG82[2]\ : NOR3C
      port map(A => \U2/un1_cnt_3\, B => \U2/un1_cnt_4\, C => 
        \U2/un1_cnt_8\, Y => \U2/un1_cnt\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I77_Y_1\ : AO1
      port map(A => \U1/N231\, B => \U1/N234\, C => 
        \U1/ADD_14x14_fast_I77_Y_0\, Y => 
        \U1/ADD_14x14_fast_I77_Y_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I20_Y\ : AO1
      port map(A => \U1/N197\, B => \U1/N201\, C => \U1/N200\, Y
         => \U1/N236\);
    
    \U0/data_ad_RNO[7]\ : NOR2A
      port map(A => \data_in_c[7]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[7]\);
    
    \U3/cnt[5]\ : DFN1C0
      port map(D => \U3/cnt_4[5]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U3/cnt[5]_net_1\);
    
    \U4/addr_RNIHVDN[2]\ : NOR2B
      port map(A => \U4/N_8_0\, B => \addr_c[2]\, Y => \U4/N_9_0\);
    
    \U1/data_all_RNO[55]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2147\, C
         => \U1/N_2148\, Y => \U1/N_692\);
    
    \U1/data_all_RNO[111]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[111]\, 
        C => \U1/N_829\, Y => \U1/N_1608\);
    
    \U1/data_all[70]\ : DFN1E0C0
      port map(D => \U1/N_175\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[70]\);
    
    \U1/pr_state_RNO[4]\ : NOR2A
      port map(A => \U1/pr_state[5]_net_1\, B => \U1/N_1084\, Y
         => \U1/pr_state_ns[3]\);
    
    \U1/data_filter_RNO[11]\ : OA1C
      port map(A => \U1/pr_state_0[5]_net_1\, B => 
        \U1/un2_data_filter[11]\, C => 
        \U1/data_filter_4_i_0_0_0[11]\, Y => \U1/N_35\);
    
    \U1/data_all[213]\ : DFN1E0C0
      port map(D => \U1/N_186\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[213]\);
    
    \data_in_pad[5]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[5]/U0/NET1\, Y => 
        \data_in_c[5]\);
    
    \U5/data_send_RNO_26[6]\ : MX2
      port map(A => \data_all[198]\, B => \data_all[206]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_441\);
    
    \U0/data_ad[11]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[11]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[11]\);
    
    \U1/data_all_RNO[213]\ : OA1B
      port map(A => \U1/N_840\, B => \U1/data_filter[5]_net_1\, C
         => \U1/data_all_3_0_0_i_0[213]\, Y => \U1/N_186\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I7_G0N\ : NOR2B
      port map(A => \data_ad[7]\, B => \U1/data_filter[7]_net_1\, 
        Y => \U1/N197\);
    
    \U2/parity_check_RNO\ : NOR3
      port map(A => \U2/parity_check_10_iv_0_3\, B => 
        \U2/parity_check_10_iv_0_2\, C => 
        \U2/parity_check_10_iv_0_4\, Y => \U2/parity_check_10_iv\);
    
    \U1/data_all[153]\ : DFN1E0C0
      port map(D => \U1/N_1799\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[153]\);
    
    \U1/pr_state_RNO_2[3]\ : NOR2A
      port map(A => \U1/N_857\, B => addr_over, Y => \U1/N_869\);
    
    \U0/ce_RNO\ : NOR2
      port map(A => \U0/pr_state[2]_net_1\, B => 
        \U0/pr_state[5]_net_1\, Y => \U0/N_138\);
    
    \U5/cnt_RNIOMCF1[4]\ : NOR3C
      port map(A => \U5/cnt[3]_net_1\, B => \U5/cnt[4]_net_1\, C
         => \U5/cnt[2]_net_1\, Y => \U5/m7_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I10_P0N\ : OR2
      port map(A => \data_ad[10]\, B => 
        \U1/data_filter[10]_net_1\, Y => \U1/N207\);
    
    \U1/data_all[83]\ : DFN1E0C0
      port map(D => \U1/N_212\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[83]\);
    
    \U3/un7_cnt_1_I_27\ : AND3
      port map(A => \U3/DWACT_FINC_E[4]\, B => \U3/cnt[8]_net_1\, 
        C => \U3/cnt[9]_net_1\, Y => \U3/N_3\);
    
    \U1/data_all[76]\ : DFN1E0C0
      port map(D => \U1/N_187\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[76]\);
    
    \U1/pr_state[2]\ : DFN1C0
      port map(D => \U1/pr_state[4]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U1/pr_state_0[2]\);
    
    \U1/data_all_RNO_1[153]\ : NOR2
      port map(A => \U1/data_filter[9]_net_1\, B => \U1/N_842\, Y
         => \U1/N_2232\);
    
    \U1/data_all_RNO[238]\ : NOR3C
      port map(A => \data_all[238]\, B => \U1/pr_state[2]_net_1\, 
        C => \U1/N_837_0\, Y => \U1/N_160\);
    
    \tx_uart_pad/U0/U0\ : IOPAD_TRI
      port map(D => \tx_uart_pad/U0/NET1\, E => 
        \tx_uart_pad/U0/NET2\, PAD => tx_uart);
    
    \U3/cnt[2]\ : DFN1C0
      port map(D => \U3/I_7\, CLK => sys_clk_c, CLR => sys_rest_c, 
        Q => \U3/cnt[2]_net_1\);
    
    \U1/cnt_daly_RNIBNTG2[5]\ : OR2A
      port map(A => \U1/cnt_daly[5]_net_1\, B => \U1/N_848\, Y
         => \U1/N_849\);
    
    \U5/data_send_RNO_24[7]\ : MX2
      port map(A => \data_all[167]\, B => \data_all[175]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_426\);
    
    \U5/data_send_RNO_18[4]\ : MX2
      port map(A => \data_all[68]\, B => \data_all[76]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_375\);
    
    \U3/data_recive_RNO_0[1]\ : NOR2A
      port map(A => \data_recive[1]\, B => send_over, Y => 
        \U3/m91_0\);
    
    \U1/cnt_daly_RNIVDVQ[8]\ : NOR2B
      port map(A => \U1/cnt_daly[8]_net_1\, B => 
        \U1/cnt_daly[3]_net_1\, Y => \U1/m24_m4_e_2\);
    
    \U1/data_all_RNO_0[9]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[9]\, Y => 
        \U1/N_1077\);
    
    \U1/data_all_RNO[141]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[141]\, Y => \U1/N_97\);
    
    \U2/parity_check_RNO_11\ : AO1A
      port map(A => \U2/N_55_i\, B => \U2/parity_check_7_sqmuxa\, 
        C => \U2/N_118\, Y => \U2/parity_check_10_iv_0_1\);
    
    \U1/data_all[107]\ : DFN1E0C0
      port map(D => \U1/N_44\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[107]\);
    
    \U1/data_all[75]\ : DFN1E0C0
      port map(D => \U1/N_185\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[75]\);
    
    \data_in_pad[4]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[4]/U0/NET1\, Y => 
        \data_in_c[4]\);
    
    \U3/cnt_RNIQUUF[11]\ : NOR2B
      port map(A => \U3/cnt[11]_net_1\, B => \U3/cnt[2]_net_1\, Y
         => \U3/m106_0\);
    
    \U1/data_all_RNO_0[226]\ : AO1C
      port map(A => \data_all[226]\, B => \U1/N_837_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m98_1_i_0\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I8_G0N\ : NOR2B
      port map(A => \data_ad[8]\, B => \U1/data_filter[8]_net_1\, 
        Y => \U1/N200\);
    
    \U1/data_all[188]\ : DFN1E0C0
      port map(D => \U1/N_417\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[188]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I31_Y\ : NOR2B
      port map(A => \U1/N186\, B => \U1/N183\, Y => \U1/N247\);
    
    \U3/cnt[4]\ : DFN1C0
      port map(D => \U3/I_12\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/cnt[4]_net_1\);
    
    \U2/cnt_RNI767T[10]\ : NOR2A
      port map(A => \U2/cnt[10]_net_1\, B => \U2/cnt[11]_net_1\, 
        Y => \U2/N_177\);
    
    \U1/data_all_RNO_0[57]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[57]\, Y => 
        \U1/N_2143\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I96_Y\ : AX1D
      port map(A => \U1/N265\, B => \U1/I68_un1_Y\, C => 
        \U1/ADD_14x14_fast_I96_Y_0\, Y => \U1/un2_data_filter[8]\);
    
    \U1/data_all_RNO_0[237]\ : AO1C
      port map(A => \data_all[237]\, B => \U1/N_837_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m69_i_0_0\);
    
    \U1/data_all_RNO[22]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/m147_0_0_i_0\, Y => \U1/N_772\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I2_G0N\ : NOR2B
      port map(A => \data_ad[2]\, B => \U1/data_filter[2]_net_1\, 
        Y => \U1/N182\);
    
    \U5/data_send_RNO_5[0]\ : MX2
      port map(A => \U5/N_507\, B => \U5/N_74\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_75\);
    
    \U2/cnt_RNIDHE91[0]\ : NOR2B
      port map(A => \U2/N_126\, B => \U2/N_168\, Y => \U2/N_174\);
    
    \U1/data_all_RNO_1[27]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_836\, 
        Y => \U1/N_2256\);
    
    \U5/data_send_RNO_16[1]\ : MX2
      port map(A => \data_all[33]\, B => \data_all[41]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_356\);
    
    \U5/data_send_RNO_8[1]\ : MX2
      port map(A => \U5/N_372\, B => \U5/N_380\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_476\);
    
    \U1/data_all_RNO_1[76]\ : NOR2
      port map(A => \U1/data_filter[12]_net_1\, B => \U1/N_833\, 
        Y => \U1/N_956\);
    
    \U5/cnt_RNIIGCF1[2]\ : NOR2B
      port map(A => \U5/N_10_0\, B => \U5/cnt[2]_net_1\, Y => 
        \U5/N_11_0\);
    
    \U1/data_all_RNO[226]\ : OA1B
      port map(A => \U1/N_837_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/m98_1_i_0\, Y => \U1/N_706\);
    
    \U1/data_all[203]\ : DFN1E0C0
      port map(D => \U1/N_75\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[203]\);
    
    \U1/cnt_daly[10]\ : DFN1E0C0
      port map(D => \U1/cnt_daly_n10\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => 
        \U1/cnt_daly[10]_net_1\);
    
    \U2/cnt_RNISS7J[1]\ : NOR3A
      port map(A => \U2/N_166\, B => \U2/cnt[6]_net_1\, C => 
        \U2/cnt[1]_net_1\, Y => \U2/tx_uart27_0_a2_2\);
    
    \U1/data_all_RNO_0[123]\ : AO1C
      port map(A => \data_all[123]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[123]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I92_Y\ : XOR3
      port map(A => \U1/data_filter[4]_net_1\, B => \data_ad[4]\, 
        C => \U1/N273\, Y => \U1/un2_data_filter[4]\);
    
    \U1/m206_i_0_o2_1\ : OR3A
      port map(A => \U1/I_7_0\, B => \U1/OVER\, C => \U1/I_9_0\, 
        Y => \U1/N_826\);
    
    \U5/data_send_RNO_19[7]\ : MX2
      port map(A => \data_all[87]\, B => \data_all[95]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_386\);
    
    \U3/un7_cnt_1_I_24\ : AND3
      port map(A => \U3/DWACT_FINC_E[0]\, B => 
        \U3/DWACT_FINC_E[2]\, C => \U3/DWACT_FINC_E[3]\, Y => 
        \U3/DWACT_FINC_E[4]\);
    
    \U1/data_all[131]\ : DFN1E0C0
      port map(D => \U1/N_78\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[131]\);
    
    \U1/data_all_RNO[189]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[189]\, Y => \U1/N_419\);
    
    \U1/data_all[13]\ : DFN1E0C0
      port map(D => \U1/N_787\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[13]\);
    
    \U3/cnt_RNIEAUG[2]\ : NOR2A
      port map(A => \U3/cnt[2]_net_1\, B => \U3/cnt[6]_net_1\, Y
         => \U3/m17_0\);
    
    \U2/idle_send_RNO_0\ : NOR2A
      port map(A => \U2/send_net_1\, B => \U2/un1_tx_uart27\, Y
         => \U2/idle_send_2_sqmuxa\);
    
    \U1/data_all[198]\ : DFN1E0C0
      port map(D => \U1/N_206\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[198]\);
    
    \U1/data_all_RNO_1[90]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_834\, 
        Y => \U1/N_2292\);
    
    \U1/data_all_RNO_1[187]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_844\, 
        Y => \U1/N_2080\);
    
    \U5/data_send_RNO_14[6]\ : MX2
      port map(A => \data_all[6]\, B => \data_all[14]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_345\);
    
    \U5/data_send_RNO[1]\ : MX2A
      port map(A => \U5/i61_mux\, B => \U5/N_69\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[1]\);
    
    \U1/data_all_RNO_0[205]\ : AO1C
      port map(A => \data_all[205]\, B => \U1/N_839_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m106_i_0_0\);
    
    \U1/data_all[88]\ : DFN1E0C0
      port map(D => \U1/N_202\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[88]\);
    
    \U2/cnt_RNI6QQV_0[10]\ : NOR3A
      port map(A => \U2/send_net_1\, B => \U2/cnt[11]_net_1\, C
         => \U2/cnt[10]_net_1\, Y => \U2/N_127\);
    
    \U1/data_all_RNO_1[5]\ : NOR2
      port map(A => \U1/data_filter[5]_net_1\, B => \U1/N_835\, Y
         => \U1/N_1087\);
    
    \U1/data_filter_RNO[9]\ : OA1C
      port map(A => \U1/pr_state_0[5]_net_1\, B => 
        \U1/un2_data_filter[9]\, C => \U1/m45_0_0_0\, Y => 
        \U1/N_46_0\);
    
    \U1/data_all_RNO[1]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1098\, C
         => \U1/N_1099\, Y => \U1/N_261\);
    
    \U1/data_all_RNO[164]\ : OA1B
      port map(A => \U1/N_838\, B => \U1/data_filter[4]_net_1\, C
         => \U1/m182_i_0_0\, Y => \U1/N_315\);
    
    \U5/data_send_RNO_28[6]\ : MX2
      port map(A => \data_all[230]\, B => \data_all[238]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_457\);
    
    \U2/parity_check_RNO_3\ : OR3
      port map(A => \U2/tx_uart36\, B => \U2/tx_uart27\, C => 
        \U2/un1_tx_uart27_6\, Y => \U2/un1_tx_uart27_1_1\);
    
    \U1/data_all_RNO[77]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m212_0_i_0\, Y => \U1/N_724\);
    
    \U2/cnt_n8\ : XA1
      port map(A => \U2/cnt_c7_net_1\, B => \U2/cnt[8]_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n8_net_1\);
    
    \U1/un14_data_all_I_7\ : AX1B
      port map(A => \addr_c[1]\, B => \addr_c[0]\, C => 
        \addr_c[2]\, Y => \U1/I_7_0\);
    
    \U4/pr_state[1]\ : DFN1C0
      port map(D => \U4/nx_state[1]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U4/pr_state[1]_net_1\);
    
    \U1/data_all_RNO_0[55]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[55]\, Y => 
        \U1/N_2147\);
    
    \U1/data_all_RNO_0[76]\ : NOR2A
      port map(A => \U1/N_833\, B => \data_all[76]\, Y => 
        \U1/N_955\);
    
    \U1/data_all[237]\ : DFN1E0C0
      port map(D => \U1/N_227\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[237]\);
    
    \U1/data_all_RNO_1[33]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_832\, Y
         => \U1/N_2218\);
    
    \U1/data_all_RNO_0[170]\ : AO1C
      port map(A => \data_all[170]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m164_i_0_0\);
    
    \U1/data_all[53]\ : DFN1E0C0
      port map(D => \U1/N_48\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[53]\);
    
    \U1/data_all_RNO_0[68]\ : NOR2A
      port map(A => \U1/N_833\, B => \data_all[68]\, Y => 
        \U1/N_971\);
    
    \U3/data_recive_RNO_0[0]\ : NOR2A
      port map(A => \data_recive[0]\, B => send_over, Y => 
        \U3/m93_0\);
    
    \data_in_pad[10]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[10]/U0/NET1\, Y => 
        \data_in_c[10]\);
    
    \U1/data_all_RNO[7]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[7]\, Y => \U1/N_248\);
    
    \U5/data_send_RNO_25[1]\ : MX2
      port map(A => \data_all[177]\, B => \data_all[185]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_428\);
    
    \U1/data_all[216]\ : DFN1E0C0
      port map(D => \U1/N_1779\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[216]\);
    
    \U3/cnt_RNI8BEO_0[11]\ : NOR3
      port map(A => \U3/cnt[4]_net_1\, B => \U3/cnt[9]_net_1\, C
         => \U3/cnt[11]_net_1\, Y => \U3/N_39\);
    
    \U3/cnt_RNI8BEO[11]\ : NOR3B
      port map(A => \U3/cnt[9]_net_1\, B => \U3/cnt[4]_net_1\, C
         => \U3/cnt[11]_net_1\, Y => \U3/N_110_mux\);
    
    \U1/data_all_RNO_0[140]\ : AO1C
      port map(A => \data_all[140]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[140]\);
    
    \U5/data_send_RNO_22[2]\ : MX2
      port map(A => \data_all[130]\, B => \data_all[138]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_405\);
    
    \U1/data_all_RNO_1[225]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_837\, Y
         => \U1/N_2164\);
    
    \U5/data_send_RNO_0[2]\ : MX2C
      port map(A => \U5/N_517\, B => \U5/N_525\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i63_mux\);
    
    \U1/data_all_RNO[87]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2135\, C
         => \U1/N_2136\, Y => \U1/N_358\);
    
    \U0/conver_ris_RNO\ : OR2B
      port map(A => \U0/conver_ris3_i_0\, B => 
        \U0/conver_ris2_net_1\, Y => \U0/conver_ris_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I78_un1_Y_0\ : NOR3C
      port map(A => \U1/N237\, B => \U1/N233\, C => \U1/N268\, Y
         => \U1/ADD_14x14_fast_I78_un1_Y_0\);
    
    \U1/data_all_RNO_0[61]\ : AO1C
      port map(A => \data_all[61]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[61]\);
    
    \U1/data_all_RNO_0[28]\ : NOR2A
      port map(A => \U1/N_836\, B => \data_all[28]\, Y => 
        \U1/N_2253\);
    
    \U1/data_all[121]\ : DFN1E0C0
      port map(D => \U1/N_382\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[121]\);
    
    \U5/cnt[2]\ : DFN1E0C0
      port map(D => \U5/cnt_n2\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \U5/cnt[2]_net_1\);
    
    \U1/data_filter[12]\ : DFN1E0C0
      port map(D => \U1/data_filter_4[12]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[12]_net_1\);
    
    \U3/cnt_RNIKFN33[0]\ : OR3C
      port map(A => \U3/m106_6\, B => \U3/m106_5\, C => 
        \U3/m106_7\, Y => \U3/un1_cnt\);
    
    \U2/cnt_RNI8PAD2_0[10]\ : NOR3C
      port map(A => \U2/N_154\, B => \U2/N_153\, C => \U2/N_178\, 
        Y => \U2/N_112\);
    
    \U1/data_all_RNO[122]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[122]\, Y => \U1/N_384\);
    
    \U2/cnt_RNI7NJ9_1[0]\ : NOR2
      port map(A => \U2/cnt[0]_net_1\, B => \U2/cnt[3]_net_1\, Y
         => \U2/N_165\);
    
    \U1/data_all_RNO[71]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/m231_i_0_0\, Y => \U1/N_177\);
    
    \U3/rx_fall\ : DFN1C0
      port map(D => rx_uart_c, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/rx_fall_net_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I62_un1_Y\ : NOR3C
      port map(A => \U1/N237\, B => \U1/N233\, C => \U1/N267\, Y
         => \U1/I62_un1_Y\);
    
    \U1/data_all[211]\ : DFN1E0C0
      port map(D => \U1/N_192\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[211]\);
    
    \U1/data_all[113]\ : DFN1E0C0
      port map(D => \U1/N_366\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[113]\);
    
    \U1/cnt_daly[2]\ : DFN1E0C0
      port map(D => \U1/N_798\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[2]_net_1\);
    
    \U2/cnt_n7\ : XA1
      port map(A => \U2/cnt_c6_net_1\, B => \U2/cnt[7]_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n7_net_1\);
    
    \U1/data_all_RNO[174]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_838\, C
         => \data_all[174]\, Y => \U1/data_all_3[174]\);
    
    \U1/data_all[82]\ : DFN1E0C0
      port map(D => \U1/N_216\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[82]\);
    
    \U1/data_all[150]\ : DFN1E0C0
      port map(D => \U1/N_751\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[150]\);
    
    \U1/data_all_RNO_0[21]\ : AO1C
      port map(A => \data_all[21]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m150_i_0_0\);
    
    \U1/data_all_RNO[49]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2155\, C
         => \U1/N_2156\, Y => \U1/N_700\);
    
    \data_in_pad[11]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[11]/U0/NET1\, Y => 
        \data_in_c[11]\);
    
    \U1/data_all[227]\ : DFN1E0C0
      port map(D => \U1/N_704\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[227]\);
    
    \U1/data_all_RNO_1[227]\ : NOR2
      port map(A => \U1/data_filter[3]_net_1\, B => \U1/N_837\, Y
         => \U1/N_2160\);
    
    \U1/data_all_RNO[154]\ : OA1B
      port map(A => \U1/N_842\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/m88_0_i_0_0\, Y => \U1/N_1800\);
    
    \U3/data_recive_RNO_3[3]\ : NOR3A
      port map(A => \U3/cnt[7]_net_1\, B => \U3/cnt[10]_net_1\, C
         => \U3/cnt[3]_net_1\, Y => \U3/m36_3\);
    
    \U1/data_all_3_0_0_i_o2_0[92]\ : OR2
      port map(A => \U1/I_5_0\, B => \addr_c[0]\, Y => \U1/N_821\);
    
    \U5/data_send_RNO_28[0]\ : MX2
      port map(A => \data_all[224]\, B => \data_all[232]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_451\);
    
    \U1/data_all_RNO_0[155]\ : AO1C
      port map(A => \data_all[155]\, B => \U1/N_842_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m83_1_i_0_0\);
    
    \U1/data_all_RNO[33]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2217\, C
         => \U1/N_2218\, Y => \U1/N_154\);
    
    \U5/data_send_RNO_3[2]\ : MX2
      port map(A => \U5/N_477\, B => \U5/N_485\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_525\);
    
    \U5/data_send_RNO_25[5]\ : MX2
      port map(A => \data_all[181]\, B => \data_all[189]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_432\);
    
    \U2/cnt_n1\ : XA1
      port map(A => \U2/cnt[1]_net_1\, B => \U2/cnt[0]_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n1_net_1\);
    
    \U1/data_all_RNO_1[68]\ : NOR2
      port map(A => \U1/data_filter[4]_net_1\, B => \U1/N_833\, Y
         => \U1/N_972\);
    
    \U1/data_all[18]\ : DFN1E0C0
      port map(D => \U1/N_1784\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[18]\);
    
    \U1/data_all[184]\ : DFN1E0C0
      port map(D => \U1/N_409\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[184]\);
    
    \U3/un7_cnt_1_I_15\ : AND2
      port map(A => \U3/cnt[3]_net_1\, B => \U3/cnt[4]_net_1\, Y
         => \U3/DWACT_FINC_E[1]\);
    
    \U2/cnt_RNI9QRS[2]\ : NOR2B
      port map(A => \U2/N_131\, B => \U2/N_172\, Y => \U2/N_178\);
    
    \U1/data_all_RNO[81]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2073\, C
         => \U1/N_1050\, Y => \U1/N_220\);
    
    \U5/data_send_RNO_11[0]\ : MX2
      port map(A => \U5/N_419\, B => \U5/N_427\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_499\);
    
    \U5/data_send_RNO_9[7]\ : MX2
      port map(A => \U5/N_394\, B => \U5/N_402\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_490\);
    
    \U3/cnt[6]\ : DFN1C0
      port map(D => \U3/cnt_4[6]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U3/cnt[6]_net_1\);
    
    \U1/data_all_RNO[25]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/m138_0_i_0_0\, Y => \U1/N_1790\);
    
    \U2/cnt_n4_tz\ : AX1C
      port map(A => \U2/cnt[3]_net_1\, B => \U2/cnt_c2_net_1\, C
         => \U2/cnt[4]_net_1\, Y => \U2/cnt_n4_tz_net_1\);
    
    \U1/data_all[0]\ : DFN1E0C0
      port map(D => \U1/N_264\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[0]\);
    
    \U5/data_send_RNO_26[5]\ : MX2
      port map(A => \data_all[197]\, B => \data_all[205]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_440\);
    
    \U1/cnt_daly_RNO_0[8]\ : OR3B
      port map(A => \U1/cnt_daly[7]_net_1\, B => 
        \U1/cnt_daly[8]_net_1\, C => \U1/N_850\, Y => \U1/N_852\);
    
    \U5/data_send_RNO_19[5]\ : MX2
      port map(A => \data_all[85]\, B => \data_all[93]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_384\);
    
    \U1/data_all_RNO[67]\ : OA1B
      port map(A => \U1/N_833\, B => \U1/data_filter[3]_net_1\, C
         => \U1/m243_i_0_0\, Y => \U1/N_169\);
    
    \U5/cnt_0[2]\ : DFN1E0C0
      port map(D => \U5/cnt_n2\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \U5/cnt_0[2]_net_1\);
    
    \U1/data_all[206]\ : DFN1E0C0
      port map(D => \U1/N_49\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[206]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I76_Y_1\ : AO1
      port map(A => \U1/N256\, B => \U1/N263\, C => 
        \U1/ADD_14x14_fast_I76_Y_0\, Y => 
        \U1/ADD_14x14_fast_I76_Y_1\);
    
    \U1/data_all_RNO_0[230]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[230]\, Y => 
        \U1/N_915\);
    
    \U1/data_all[232]\ : DFN1E0C0
      port map(D => \U1/N_221\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[232]\);
    
    \U1/data_all_RNO[204]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[204]\, Y => \U1/N_100\);
    
    \U2/cnt_c4\ : NOR3C
      port map(A => \U2/cnt[3]_net_1\, B => \U2/cnt_c2_net_1\, C
         => \U2/cnt[4]_net_1\, Y => \U2/cnt_c4_net_1\);
    
    \U1/data_all[79]\ : DFN1E0C0
      port map(D => \U1/data_all_3[79]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[79]\);
    
    \U2/cnt_RNIVV7J[8]\ : NOR3C
      port map(A => \U2/cnt[7]_net_1\, B => \U2/cnt[8]_net_1\, C
         => \U2/tx_uart36_5\, Y => \U2/tx_uart36_8\);
    
    \U1/data_all[58]\ : DFN1E0C0
      port map(D => \U1/N_686\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[58]\);
    
    \U1/ad_once_over_RNO\ : NOR3
      port map(A => \U1/pr_state_0[7]_net_1\, B => 
        \U1/pr_state[4]_net_1\, C => \U1/pr_state[2]_net_1\, Y
         => \U1/N_1092\);
    
    \U1/data_all[81]\ : DFN1E0C0
      port map(D => \U1/N_220\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[81]\);
    
    \U1/data_all[34]\ : DFN1E0C0
      port map(D => \U1/N_1807\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[34]\);
    
    \U5/data_send_RNO_10[6]\ : MX2
      port map(A => \U5/N_409\, B => \U5/N_417\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_497\);
    
    \U5/data_send_RNO_3[3]\ : MX2
      port map(A => \U5/N_478\, B => \U5/N_486\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_526\);
    
    \U4/nx_state_RNO[0]\ : AXOI5
      port map(A => \U4/N_11_0\, B => \U4/pr_state[0]_net_1\, C
         => \U4/pr_state[1]_net_1\, Y => 
        \U4/nx_state_RNO[0]_net_1\);
    
    \U2/tx_uart\ : DFN1E0P0
      port map(D => \U2/tx_uart_11\, CLK => sys_clk_c, PRE => 
        sys_rest_c, E => \U2/tx_uart_11_sqmuxa\, Q => tx_uart_c);
    
    \U1/data_all[87]\ : DFN1E0C0
      port map(D => \U1/N_358\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[87]\);
    
    \U2/cnt_RNI7DUF2[10]\ : NOR3C
      port map(A => \U2/N_169\, B => \U2/N_127\, C => \U2/N_180\, 
        Y => \U2/parity_check_3_sqmuxa\);
    
    \tx_uart_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => tx_uart_c, E => \VCC\, DOUT => 
        \tx_uart_pad/U0/NET1\, EOUT => \tx_uart_pad/U0/NET2\);
    
    \U5/data_send_RNO_2[1]\ : MX2
      port map(A => \U5/N_460\, B => \U5/N_468\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_516\);
    
    \U1/data_all_RNO[59]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2139\, C
         => \U1/N_2140\, Y => \U1/N_680\);
    
    \U1/data_all[30]\ : DFN1E0C0
      port map(D => \U1/data_all_3[30]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[30]\);
    
    \U1/data_all[201]\ : DFN1E0C0
      port map(D => \U1/N_2041\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[201]\);
    
    \U1/data_all[103]\ : DFN1E0C0
      port map(D => \U1/N_52\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[103]\);
    
    \U1/data_all_RNO[98]\ : OA1B
      port map(A => \U1/N_829\, B => \U1/data_filter[2]_net_1\, C
         => \U1/data_all_3_i_0_0_0[98]\, Y => \U1/N_1613\);
    
    \U1/data_all[194]\ : DFN1E0C0
      port map(D => \U1/N_93\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[194]\);
    
    \U1/data_all_RNO[139]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[11]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[139]\, Y => \U1/N_1837\);
    
    \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_1[63]\ : OR2A
      port map(A => \U1/I_5_0\, B => \U1/I_9_0\, Y => \U1/N_820\);
    
    \U1/data_all[12]\ : DFN1E0C0
      port map(D => \U1/N_239\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[12]\);
    
    \U1/cnt_daly_RNIFDGQ[11]\ : NOR2A
      port map(A => \U1/cnt_daly[9]_net_1\, B => 
        \U1/cnt_daly[11]_net_1\, Y => \U1/m61_0_i_a3_1_1\);
    
    \data_in_pad[7]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[7]/U0/NET1\, Y => 
        \data_in_c[7]\);
    
    \U2/cnt_RNI0ISQ4[8]\ : AO1
      port map(A => \U2/tx_uart37_8\, B => \U2/tx_uart37_7\, C
         => \U2/tx_uart38\, Y => \U2/un1_tx_uart27_6\);
    
    \U0/data_ad_RNO[11]\ : NOR2A
      port map(A => \data_in_c[11]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[11]\);
    
    \U5/data_send_RNO_24[0]\ : MX2
      port map(A => \data_all[160]\, B => \data_all[168]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_419\);
    
    \U1/data_all_RNO_0[156]\ : AO1C
      port map(A => \data_all[156]\, B => \U1/N_842\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m82_1_i_i_0\);
    
    \U1/data_all_RNO[61]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[61]\, Y => \U1/N_356\);
    
    \U1/data_all[138]\ : DFN1E0C0
      port map(D => \U1/N_101\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[138]\);
    
    \U1/cnt_daly[4]\ : DFN1E0C0
      port map(D => \U1/N_802\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[4]_net_1\);
    
    \U3/cnt_4[6]\ : XA1
      port map(A => \U3/N_7\, B => \U3/cnt[6]_net_1\, C => 
        \U3/recive_net_1\, Y => \U3/cnt_4[6]_net_1\);
    
    \U1/data_all_RNO_0[152]\ : AO1C
      port map(A => \data_all[152]\, B => \U1/N_842\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m92_1_i_0_0\);
    
    \U1/data_all[36]\ : DFN1E0C0
      port map(D => \U1/N_1809\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[36]\);
    
    \U2/parity_check_RNO_1\ : AO1A
      port map(A => \U2/N_68_i\, B => \U2/parity_check_3_sqmuxa\, 
        C => \U2/N_120\, Y => \U2/parity_check_10_iv_0_3\);
    
    \U0/pr_state[2]\ : DFN1C0
      port map(D => \U0/pr_state_RNO[2]_net_1\, CLK => sys_clk_c, 
        CLR => sys_rest_c, Q => \U0/pr_state[2]_net_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I1_G0N\ : NOR2B
      port map(A => \data_ad[1]\, B => \U1/data_filter[1]_net_1\, 
        Y => \U1/N179\);
    
    \U1/data_all_RNO_0[12]\ : AO1C
      port map(A => \data_all[12]\, B => \U1/N_835_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[12]\);
    
    \U1/data_all_RNO[199]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/m124_0_i_0\, Y => \U1/N_85\);
    
    \U1/data_all_3_0_a2_i_0_o2_0_0[239]\ : OR2
      port map(A => \U1/m146_i_0_o2_1\, B => \U1/N_818\, Y => 
        \U1/N_837_0\);
    
    \U2/cnt_RNI8PAD2[10]\ : NOR3C
      port map(A => \U2/N_154\, B => \U2/N_153\, C => \U2/N_196\, 
        Y => \U2/N_114\);
    
    \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_0_0[63]\ : OR2
      port map(A => 
        \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_0[63]_net_1\, B => 
        \U1/N_817\, Y => \U1/N_831_0\);
    
    \U1/data_all[222]\ : DFN1E0C0
      port map(D => \U1/N_1781\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[222]\);
    
    \U1/data_all[52]\ : DFN1E0C0
      port map(D => \U1/N_694\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[52]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I16_Y\ : AO1
      port map(A => \U1/N203\, B => \U1/N207\, C => \U1/N206\, Y
         => \U1/N232\);
    
    \U5/data_send_RNO_1[0]\ : MX2A
      port map(A => \U5/N_537\, B => \U5/N_75\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_76\);
    
    \U5/data_send_RNO_21[3]\ : MX2
      port map(A => \data_all[115]\, B => \data_all[123]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_398\);
    
    \U3/data_recive[5]\ : DFN1C0
      port map(D => \U3/data_recive_12[5]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[5]\);
    
    \U1/data_all_RNO[32]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/m298_i_0_0\, Y => \U1/N_1806\);
    
    \U1/data_all[35]\ : DFN1E0C0
      port map(D => \U1/N_1808\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[35]\);
    
    \U5/data_send_RNO_19[4]\ : MX2
      port map(A => \data_all[84]\, B => \data_all[92]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_383\);
    
    \U5/data_send_RNO_12[7]\ : MX2
      port map(A => \U5/N_442\, B => \U5/N_450\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_514\);
    
    \U2/cnt_RNISS7J_2[1]\ : NOR2B
      port map(A => \U2/N_128\, B => \U2/N_164\, Y => \U2/N_172\);
    
    \U5/data_send_RNO_25[2]\ : MX2
      port map(A => \data_all[178]\, B => \data_all[186]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_429\);
    
    \U1/data_all[1]\ : DFN1E0C0
      port map(D => \U1/N_261\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[1]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I12_Y\ : NOR3C
      port map(A => \U1/data_filter[11]_net_1\, B => 
        \data_ad[11]\, C => \U1/data_filter[12]_net_1\, Y => 
        \U1/N227\);
    
    \U1/data_all_RNO_1[233]\ : NOR2
      port map(A => \U1/data_filter[9]_net_1\, B => \U1/N_837_0\, 
        Y => \U1/N_912\);
    
    \U1/data_all_RNO[116]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[116]\, Y => \U1/N_372\);
    
    \U5/data_send_RNO_17[2]\ : MX2
      port map(A => \data_all[50]\, B => \data_all[58]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_365\);
    
    \U1/data_all_RNO_0[218]\ : AO1C
      port map(A => \data_all[218]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[218]\);
    
    \U1/data_all[11]\ : DFN1E0C0
      port map(D => \U1/N_241\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[11]\);
    
    \U3/data_recive_RNO_4[0]\ : NOR3B
      port map(A => \U3/cnt[6]_net_1\, B => \U3/cnt[2]_net_1\, C
         => \U3/cnt[3]_net_1\, Y => \U3/m62_4\);
    
    \U1/data_all[17]\ : DFN1E0C0
      port map(D => \U1/N_1783\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[17]\);
    
    \U5/data_send_RNO_22[3]\ : MX2
      port map(A => \data_all[131]\, B => \data_all[139]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_406\);
    
    \U5/data_send_RNO_6[3]\ : MX2
      port map(A => \U5/N_342\, B => \U5/N_350\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_462\);
    
    \U4/addr[2]\ : DFN1E0C0
      port map(D => \U4/addr_n2\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U4/N_7_0\, Q => \addr_c[2]\);
    
    \U1/data_all_RNO[46]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_832\, C
         => \data_all[46]\, Y => \U1/data_all_3[46]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I77_Y_0\ : MAJ3
      port map(A => \U1/data_filter[11]_net_1\, B => 
        \data_ad[11]\, C => \U1/N206\, Y => 
        \U1/ADD_14x14_fast_I77_Y_0\);
    
    \U1/data_all[128]\ : DFN1E0C0
      port map(D => \U1/N_1835\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[128]\);
    
    \U1/pr_state[7]\ : DFN1P0
      port map(D => \U1/pr_state_RNICDI39[1]_net_1\, CLK => 
        sys_clk_c, PRE => sys_rest_c, Q => \U1/pr_state[7]_net_1\);
    
    \U5/data_send_RNO_9[4]\ : MX2
      port map(A => \U5/N_391\, B => \U5/N_399\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_487\);
    
    \U1/data_all[110]\ : DFN1E0C0
      port map(D => \U1/N_1609\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[110]\);
    
    \U1/data_all_RNO[168]\ : OA1B
      port map(A => \U1/N_838\, B => \U1/data_filter[8]_net_1\, C
         => \U1/m170_i_0_0\, Y => \U1/N_323\);
    
    \U2/cnt_c6\ : NOR3C
      port map(A => \U2/cnt[5]_net_1\, B => \U2/cnt_c4_net_1\, C
         => \U2/cnt[6]_net_1\, Y => \U2/cnt_c6_net_1\);
    
    \U1/data_all_RNO[125]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[125]\, Y => \U1/N_390\);
    
    \U0/sts_ris_RNO\ : OR2A
      port map(A => \U0/sts_ris3_net_1\, B => \U0/sts_ris2_net_1\, 
        Y => \U0/sts_ris_2\);
    
    \U1/data_all_RNO_1[186]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_844\, 
        Y => \U1/N_2082\);
    
    \U1/data_all_RNO_0[135]\ : AO1C
      port map(A => \data_all[135]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m202_0_i_0\);
    
    \U5/data_send_RNO_17[1]\ : MX2
      port map(A => \data_all[49]\, B => \data_all[57]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_364\);
    
    \U1/data_all_RNO[206]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[206]\, 
        C => \U1/N_839\, Y => \U1/N_49\);
    
    \U1/data_all[176]\ : DFN1E0C0
      port map(D => \U1/N_393\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[176]\);
    
    \U5/pr_state_RNI4CS81[1]\ : XA1
      port map(A => \U5/cnt_0[2]_net_1\, B => \U5/N_10_0\, C => 
        \U5/pr_state[1]_net_1\, Y => \U5/cnt_n2\);
    
    \U1/data_all[51]\ : DFN1E0C0
      port map(D => \U1/N_696\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[51]\);
    
    \U1/receive_on\ : DFN1E1C0
      port map(D => addr_over_i, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_260\, Q => receive_on);
    
    \U2/cnt_RNI7DUF2[1]\ : NOR3C
      port map(A => \U2/N_171\, B => 
        \U2/un1_tx_uart27_3_0_a2_3_1\, C => \U2/N_174\, Y => 
        \U2/parity_check_5_sqmuxa\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I64_un1_Y\ : NOR2B
      port map(A => \U1/N262\, B => \U1/N269\, Y => 
        \U1/I64_un1_Y\);
    
    \U1/data_all_3_i_o3_0_o2_0_o2[143]\ : OR2
      port map(A => \U1/m103_i_o2_0_o2_0_net_1\, B => \U1/N_817\, 
        Y => \U1/N_841\);
    
    \U1/data_all[57]\ : DFN1E0C0
      port map(D => \U1/N_688\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[57]\);
    
    \U0/data_ad[5]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[5]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[5]\);
    
    \U1/data_all_RNO_0[214]\ : AO1C
      port map(A => \data_all[214]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[214]\);
    
    \U0/data_ad[3]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[3]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[3]\);
    
    \U3/data_recive_RNO_1[4]\ : NOR3C
      port map(A => \U3/m53_3\, B => \U3/m53_2\, C => 
        \U3/N_120_mux\, Y => \U3/data_recive27\);
    
    \U1/receive_flag_RNO_0\ : NOR2A
      port map(A => \data_recive[0]\, B => 
        \U1/cnt_receive_over_net_1\, Y => \U1/m112_i_0_a3_0\);
    
    \U1/data_all_RNO[146]\ : OA1B
      port map(A => \U1/N_842\, B => \U1/data_filter[2]_net_1\, C
         => \U1/m112_1_i_0_0\, Y => \U1/N_1796\);
    
    \U3/cnt[10]\ : DFN1C0
      port map(D => \U3/I_28\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/cnt[10]_net_1\);
    
    \U2/cnt_RNI5MRS[0]\ : NOR3C
      port map(A => \U2/N_166\, B => \U2/N_124\, C => 
        \U2/tx_uart35_0_a2_0_0\, Y => \U2/tx_uart35_0_a2_0_1\);
    
    \U1/data_all_RNO[212]\ : OA1B
      port map(A => \U1/N_840\, B => \U1/data_filter[4]_net_1\, C
         => \U1/data_all_3_0_0_i_0[212]\, Y => \U1/N_190\);
    
    \U5/data_send_RNO_20[7]\ : MX2
      port map(A => \data_all[103]\, B => \data_all[111]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_394\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I4_G0N\ : NOR2B
      port map(A => \data_ad[4]\, B => \U1/data_filter[4]_net_1\, 
        Y => \U1/N188\);
    
    \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_0[63]\ : OR3A
      port map(A => \U1/I_5_0\, B => \U1/I_9_0\, C => \addr_c[0]\, 
        Y => \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_0[63]_net_1\);
    
    \U5/data_send_RNO_13[2]\ : NOR2A
      port map(A => \U5/N_453\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_60_0\);
    
    \U1/data_all_RNO_0[60]\ : AO1C
      port map(A => \data_all[60]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[60]\);
    
    \U1/un14_data_all_I_9\ : XNOR2
      port map(A => \U1/N_3\, B => \addr_c[3]\, Y => \U1/I_9_0\);
    
    \U3/cnt[0]\ : DFN1C0
      port map(D => \U3/cnt_4[0]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/cnt[0]_net_1\);
    
    \U1/data_all_RNO_0[6]\ : AO1C
      port map(A => \data_all[6]\, B => \U1/N_835_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[6]\);
    
    \U1/data_filter[10]\ : DFN1E0C0
      port map(D => \U1/N_37\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[10]_net_1\);
    
    \U1/data_all_RNO[56]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[56]\, Y => \U1/N_690\);
    
    \U3/data_recive_RNO_2[7]\ : NOR2A
      port map(A => \U3/m22_0\, B => \U3/cnt[3]_net_1\, Y => 
        \U3/m22_2\);
    
    \U1/data_all_RNO[113]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[1]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[113]\, Y => \U1/N_366\);
    
    \U1/data_all_RNO[70]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/m234_i_0_0\, Y => \U1/N_175\);
    
    \U1/data_all[63]\ : DFN1E0C0
      port map(D => \U1/N_91\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[63]\);
    
    \U1/data_all_RNO[178]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[178]\, Y => \U1/N_397\);
    
    \U1/data_all_RNO[110]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[110]\, 
        C => \U1/N_829_0\, Y => \U1/N_1609\);
    
    \U1/data_all[7]\ : DFN1E0C0
      port map(D => \U1/N_248\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[7]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I90_Y\ : XOR3
      port map(A => \U1/data_filter[2]_net_1\, B => \data_ad[2]\, 
        C => \U1/N250\, Y => \U1/un2_data_filter[2]\);
    
    \U4/addr_over\ : DFN1E0C0
      port map(D => \U4/pr_state[1]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U4/pr_state[0]_net_1\, Q => 
        addr_over);
    
    \U3/data_recive_RNO[3]\ : MX2
      port map(A => \U3/m87_0\, B => rx_uart_c, S => 
        \U3/data_recive26\, Y => \U3/data_recive_12[3]\);
    
    \U2/cnt_n11\ : AX1C
      port map(A => \U2/cnt_c9_net_1\, B => \U2/cnt_24_0_net_1\, 
        C => \U2/N_152\, Y => \U2/cnt_n11_net_1\);
    
    \U1/data_all_RNO_0[20]\ : NOR2A
      port map(A => \U1/N_836\, B => \data_all[20]\, Y => 
        \U1/N_2269\);
    
    \U1/data_all_RNO_0[183]\ : AO1C
      port map(A => \data_all[183]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[183]\);
    
    \U5/data_send_RNO_19[3]\ : MX2
      port map(A => \data_all[83]\, B => \data_all[91]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_382\);
    
    \U2/cnt_RNIDTJ9_0[2]\ : NOR2A
      port map(A => \U2/cnt[2]_net_1\, B => \U2/cnt[7]_net_1\, Y
         => \U2/N_131\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I54_Y\ : AO1
      port map(A => \U1/N247\, B => \U1/N250\, C => \U1/N246\, Y
         => \U1/N273\);
    
    \U1/data_all_RNO_0[225]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[225]\, Y => 
        \U1/N_2163\);
    
    \U5/data_send_RNO_6[5]\ : MX2
      port map(A => \U5/N_344\, B => \U5/N_352\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_464\);
    
    \U5/data_send_RNO_1[7]\ : MX2A
      port map(A => \U5/N_530\, B => \U5/N_26_0\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_27_0\);
    
    \U3/recive\ : DFN1E1C0
      port map(D => \U3/un1_cnt\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U3/un2_cnt\, Q => \U3/recive_net_1\);
    
    \U5/data_send_RNO_5[2]\ : MX2
      port map(A => \U5/N_509\, B => \U5/N_60_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_61_0\);
    
    \U3/un7_cnt_1_I_21\ : AND2
      port map(A => \U3/cnt[6]_net_1\, B => \U3/cnt[7]_net_1\, Y
         => \U3/DWACT_FINC_E[3]\);
    
    \U1/data_all_RNO_0[139]\ : AO1C
      port map(A => \data_all[139]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[139]\);
    
    \U1/data_all_RNO[158]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_842_0\, C
         => \data_all[158]\, Y => \U1/data_all_3[158]\);
    
    \U5/data_send_RNO_24[1]\ : MX2
      port map(A => \data_all[161]\, B => \data_all[169]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_420\);
    
    \U2/cnt_c9\ : NOR2B
      port map(A => \U2/cnt_c8_net_1\, B => \U2/cnt[9]_net_1\, Y
         => \U2/cnt_c9_net_1\);
    
    \U1/data_all_RNO_0[144]\ : AO1C
      port map(A => \data_all[144]\, B => \U1/N_842\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m118_0_i_1_0\);
    
    \U1/data_all_RNO_0[136]\ : AO1C
      port map(A => \data_all[136]\, B => \U1/N_841_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m199_0_i_0\);
    
    \U2/idle_send\ : DFN1E0C0
      port map(D => \U2/idle_send_0_sqmuxa\, CLK => sys_clk_c, 
        CLR => sys_rest_c, E => \U2/idle_send_2_sqmuxa\, Q => 
        \U2/idle_send_net_1\);
    
    \U1/data_all_RNO_0[187]\ : NOR2A
      port map(A => \U1/N_844\, B => \data_all[187]\, Y => 
        \U1/N_2079\);
    
    \U1/data_all[100]\ : DFN1E0C0
      port map(D => \U1/N_58\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[100]\);
    
    \U5/data_send_RNO_27[5]\ : MX2
      port map(A => \data_all[213]\, B => \data_all[221]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_448\);
    
    \U0/data_ad_RNO[0]\ : NOR2A
      port map(A => \data_in_c[0]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[0]\);
    
    \U1/data_all_RNO_0[132]\ : AO1C
      port map(A => \data_all[132]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[132]\);
    
    \U1/data_all_RNO[18]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/m159_0_i_0_0\, Y => \U1/N_1784\);
    
    \U1/data_all[230]\ : DFN1E0C0
      port map(D => \U1/N_219\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[230]\);
    
    \U1/data_all[134]\ : DFN1E0C0
      port map(D => \U1/N_82\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[134]\);
    
    \U0/cnt_rc[1]\ : DFN1E0C0
      port map(D => \U0/cnt_rc_n1_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U0/N_135\, Q => 
        \U0/cnt_rc[1]_net_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I32_Y\ : AO1
      port map(A => \U1/N179\, B => \U1/N183\, C => \U1/N182\, Y
         => \U1/N248\);
    
    \U1/data_all_RNO[80]\ : OA1B
      port map(A => \U1/N_834_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[80]\, Y => \U1/N_224\);
    
    \U2/cnt[9]\ : DFN1C0
      port map(D => \U2/cnt_n9_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[9]_net_1\);
    
    \U1/cnt_daly_RNO[7]\ : XA1C
      port map(A => \U1/cnt_daly[7]_net_1\, B => \U1/N_850\, C
         => \U1/pr_state[7]_net_1\, Y => \U1/N_808\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I78_Y_1\ : AO1
      port map(A => \U1/ADD_14x14_fast_I78_un1_Y_0\, B => 
        \U1/N275\, C => \U1/ADD_14x14_fast_I78_Y_0\, Y => 
        \U1/ADD_14x14_fast_I78_Y_1\);
    
    \U1/data_all[179]\ : DFN1E0C0
      port map(D => \U1/N_399\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[179]\);
    
    \U4/pr_state[0]\ : DFN1C0
      port map(D => \U4/nx_state[0]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U4/pr_state[0]_net_1\);
    
    \U1/data_all_RNO[102]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[102]\, Y => \U1/N_54\);
    
    \U5/data_send_RNO_16[7]\ : MX2
      port map(A => \data_all[39]\, B => \data_all[47]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_362\);
    
    \U1/data_all_RNO_0[138]\ : NOR2A
      port map(A => \U1/N_841\, B => \data_all[138]\, Y => 
        \U1/N_947\);
    
    \U3/un7_cnt_1_I_31\ : AND3
      port map(A => \U3/DWACT_FINC_E[6]\, B => \U3/cnt[9]_net_1\, 
        C => \U3/cnt[10]_net_1\, Y => \U3/N_2\);
    
    \U5/data_send[5]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[5]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[5]\);
    
    \U2/parity_check_RNO_0\ : OA1A
      port map(A => \U2/un1_tx_uart27\, B => 
        \U2/un1_tx_uart27_1_1\, C => \U2/send_net_1\, Y => 
        \U2/parity_check_0_sqmuxa\);
    
    \U1/data_all_RNO[143]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[143]\, 
        C => \U1/N_841_0\, Y => \U1/N_17\);
    
    \U5/pr_state_RNO[0]\ : AOI1
      port map(A => \U5/N_138_mux\, B => \U5/pr_state[1]_net_1\, 
        C => \U5/pr_state_ns_0_i_0[0]\, Y => \U5/N_6\);
    
    \U1/data_all_RNO_0[200]\ : AO1C
      port map(A => \data_all[200]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m121_0_0_i_0\);
    
    \U1/data_all_RNO[140]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[140]\, Y => \U1/N_94\);
    
    \U1/cnt_daly[3]\ : DFN1E0C0
      port map(D => \U1/N_800\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[3]_net_1\);
    
    \U1/data_all_RNO[127]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[127]\, 
        C => \U1/N_830_0\, Y => \U1/N_70\);
    
    \U1/data_all_RNO[35]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/m289_i_0_0\, Y => \U1/N_1808\);
    
    \U3/rx_fall2\ : DFN1C0
      port map(D => \U3/rx_fall1_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U3/rx_fall2_net_1\);
    
    \U1/data_all[215]\ : DFN1E0C0
      port map(D => \U1/N_178\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[215]\);
    
    \U1/data_all_RNO[0]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[0]\, Y => \U1/N_264\);
    
    \U5/data_send_RNO_20[5]\ : MX2
      port map(A => \data_all[101]\, B => \data_all[109]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_392\);
    
    \U1/pr_state_RNI37MS[0]\ : NOR2
      port map(A => \U1/pr_state[0]_net_1\, B => 
        \U1/pr_state[7]_net_1\, Y => \U1/N_1090\);
    
    \U1/data_all[147]\ : DFN1E0C0
      port map(D => \U1/N_122\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[147]\);
    
    \U1/data_all_RNO_0[87]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[87]\, Y => 
        \U1/N_2135\);
    
    \U1/data_all_RNO[29]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m125_0_0_i_0\, Y => \U1/N_763\);
    
    \U4/nx_state_RNO_0[1]\ : NOR3B
      port map(A => \U4/N_11_0\, B => \U4/pr_state[0]_net_1\, C
         => \U4/pr_state[1]_net_1\, Y => 
        \U4/nx_state_RNO_0[1]_net_1\);
    
    \U3/cnt[1]\ : DFN1C0
      port map(D => \U3/I_5\, CLK => sys_clk_c, CLR => sys_rest_c, 
        Q => \U3/cnt[1]_net_1\);
    
    \U2/cnt_RNIGILQ4[10]\ : OR2
      port map(A => \U2/tx_uart36\, B => \U2/N_112\, Y => 
        \U2/un1_tx_uart27_1_0\);
    
    \U1/pr_state[3]\ : DFN1C0
      port map(D => \U1/pr_state_RNO[3]_net_1\, CLK => sys_clk_c, 
        CLR => sys_rest_c, Q => \U1/pr_state[3]_net_1\);
    
    \U1/data_all[167]\ : DFN1E0C0
      port map(D => \U1/N_321\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[167]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I3_P0N\ : OR2
      port map(A => \data_ad[3]\, B => \U1/data_filter[3]_net_1\, 
        Y => \U1/N186\);
    
    \U1/data_all_RNO_0[150]\ : AO1C
      port map(A => \data_all[150]\, B => \U1/N_842_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m98_0_i_i_0\);
    
    \U1/data_all_3_i_o3_0_o2_0_o2_0_0[143]\ : OR2
      port map(A => \U1/m103_i_o2_0_o2_0_net_1\, B => \U1/N_817\, 
        Y => \U1/N_841_0\);
    
    \U4/conver_ris2\ : DFN1C0
      port map(D => \U4/conver_ris1_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U4/conver_ris2_net_1\);
    
    \U1/m302_0_i_o2\ : OR2
      port map(A => \U1/m302_0_i_o2_0_net_1\, B => \U1/N_817\, Y
         => \U1/N_835\);
    
    \U4/pr_state_RNI876C1[1]\ : NOR2
      port map(A => \U4/N_11_0\, B => \U4/pr_state[1]_net_1\, Y
         => \U4/N_25\);
    
    \U1/data_all_RNO[93]\ : OA1B
      port map(A => \U1/N_834_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[93]\, Y => \U1/N_1776\);
    
    \U1/data_all[220]\ : DFN1E0C0
      port map(D => \U1/N_166\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[220]\);
    
    \U1/data_all[124]\ : DFN1E0C0
      port map(D => \U1/N_388\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[124]\);
    
    \U0/data_ad_RNO[8]\ : NOR2A
      port map(A => \data_in_c[8]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[8]\);
    
    \U2/cnt[8]\ : DFN1C0
      port map(D => \U2/cnt_n8_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[8]_net_1\);
    
    \U1/cnt_RNI6SD3[2]\ : OR3A
      port map(A => \U1/cnt[2]_net_1\, B => \U1/cnt[0]_net_1\, C
         => \U1/cnt[1]_net_1\, Y => \U1/N_1084\);
    
    \U1/data_all[24]\ : DFN1E0C0
      port map(D => \U1/N_1789\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[24]\);
    
    \U1/data_all[39]\ : DFN1E0C0
      port map(D => \U1/N_1812\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[39]\);
    
    \U1/data_all_RNO[60]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[60]\, Y => \U1/N_31\);
    
    \U1/data_all_RNO[218]\ : OA1B
      port map(A => \U1/N_840_0\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[218]\, Y => \U1/N_1778\);
    
    \U1/data_all[68]\ : DFN1E0C0
      port map(D => \U1/N_171\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[68]\);
    
    \U0/pr_state_RNO[0]\ : NOR2
      port map(A => \U0/N_143\, B => \U0/pr_state_ns[1]\, Y => 
        \U0/pr_state_RNO_0[0]_net_1\);
    
    \U3/data_recive_RNO[1]\ : MX2
      port map(A => \U3/m91_0\, B => rx_uart_c, S => 
        \U3/data_recive24\, Y => \U3/data_recive_12[1]\);
    
    \U1/data_all_RNO_0[195]\ : AO1C
      port map(A => \data_all[195]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m136_i_0_0\);
    
    \U1/data_all_RNO[161]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[1]_net_1\, 
        C => \U1/m188_i_0_0\, Y => \U1/N_1815\);
    
    \U1/data_filter_RNO[3]\ : OA1C
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/un2_data_filter[3]\, C => 
        \U1/data_filter_4_i_0_0_0[3]\, Y => \U1/N_1421\);
    
    \U1/data_all[20]\ : DFN1E0C0
      port map(D => \U1/N_1786\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[20]\);
    
    \U1/cnt_daly[1]\ : DFN1E0C0
      port map(D => \U1/N_796\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[1]_net_1\);
    
    \U3/data_recive_RNO_0[5]\ : NOR2A
      port map(A => \data_recive[5]\, B => send_over, Y => 
        \U3/m83_0\);
    
    \U1/m107_e_1\ : NOR2A
      port map(A => \data_recive[6]\, B => \data_recive[5]\, Y
         => \U1/m107_e_1_net_1\);
    
    \U0/rc_RNO\ : NOR2
      port map(A => \U0/N_144\, B => \U0/pr_state[0]_net_1\, Y
         => \U0/N_136\);
    
    \U5/data_send_RNO_11[2]\ : MX2
      port map(A => \U5/N_421\, B => \U5/N_429\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_501\);
    
    \sys_rest_pad/U0/U0\ : IOPAD_IN
      port map(PAD => sys_rest, Y => \sys_rest_pad/U0/NET1\);
    
    \data_in_pad[1]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[1]/U0/NET1\, Y => 
        \data_in_c[1]\);
    
    \U5/data_send_RNO_3[4]\ : MX2
      port map(A => \U5/N_479\, B => \U5/N_487\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_527\);
    
    \U1/data_all_RNO_0[16]\ : AO1C
      port map(A => \data_all[16]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m163_0_i_0_0\);
    
    \U4/addr_RNO[1]\ : XA1
      port map(A => \addr_c_0[0]\, B => \addr_c[1]\, C => 
        \U4/pr_state[0]_net_1\, Y => \U4/addr_n1\);
    
    \U1/cnt_daly_RNO_1[10]\ : NOR3C
      port map(A => \U1/cnt_daly[4]_net_1\, B => 
        \U1/cnt_daly[3]_net_1\, C => \U1/m22_m4_0_a2_2\, Y => 
        \U1/m22_m4_0_a2_4\);
    
    \U1/vld_whole_RNO\ : NOR2
      port map(A => \U1/pr_state[3]_net_1\, B => 
        \U1/pr_state[7]_net_1\, Y => \U1/N_1093\);
    
    \U1/data_all_RNO_0[85]\ : AO1C
      port map(A => \data_all[85]\, B => \U1/N_834_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[85]\);
    
    \U1/data_all[5]\ : DFN1E0C0
      port map(D => \U1/N_253\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[5]\);
    
    \U0/data_ad[7]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[7]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[7]\);
    
    \U1/data_all_RNO_0[19]\ : AO1C
      port map(A => \data_all[19]\, B => \U1/N_836\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m156_0_i_0_0\);
    
    \U1/data_all[26]\ : DFN1E0C0
      port map(D => \U1/N_1791\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[26]\);
    
    \U1/data_all_RNO_1[43]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_832\, 
        Y => \U1/N_2198\);
    
    \U1/data_all[205]\ : DFN1E0C0
      port map(D => \U1/N_213\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[205]\);
    
    \U5/data_send_RNO_22[5]\ : MX2
      port map(A => \data_all[133]\, B => \data_all[141]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_408\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I24_Y\ : AO1
      port map(A => \U1/N191\, B => \U1/N195\, C => \U1/N194\, Y
         => \U1/N240\);
    
    \U2/cnt_RNIPP7J[4]\ : NOR3C
      port map(A => \U2/cnt[5]_net_1\, B => \U2/cnt[4]_net_1\, C
         => \U2/tx_uart37_3\, Y => \U2/tx_uart37_6_0\);
    
    \U5/data_send_RNO_9[5]\ : MX2
      port map(A => \U5/N_392\, B => \U5/N_400\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_488\);
    
    \U0/cnt_rclde_i_a4\ : NOR2
      port map(A => \U0/pr_state[0]_net_1\, B => 
        \U0/pr_state[4]_net_1\, Y => \U0/N_135\);
    
    \data_in_pad[9]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(9), Y => \data_in_pad[9]/U0/NET1\);
    
    \U1/data_all_RNO_1[59]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_831\, 
        Y => \U1/N_2140\);
    
    \U1/data_all[43]\ : DFN1E0C0
      port map(D => \U1/N_284\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[43]\);
    
    \U5/data_send_RNO_3[0]\ : MX2
      port map(A => \U5/N_475\, B => \U5/N_483\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_523\);
    
    \U5/data_send_RNO[2]\ : MX2A
      port map(A => \U5/i63_mux\, B => \U5/N_62_0\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[2]\);
    
    \U4/addr_RNI62K31[3]\ : NOR2B
      port map(A => \U4/N_10_0\, B => ad_once_over, Y => 
        \U4/N_11_0\);
    
    \U3/data_recive[1]\ : DFN1C0
      port map(D => \U3/data_recive_12[1]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[1]\);
    
    \U1/data_all_RNO[8]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[8]\, Y => \U1/N_246\);
    
    \U1/data_all[62]\ : DFN1E0C0
      port map(D => \U1/N_1422\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[62]\);
    
    \U1/data_all_RNO[171]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[11]_net_1\, 
        C => \U1/m161_i_0_0\, Y => \U1/N_329\);
    
    \U1/data_all[25]\ : DFN1E0C0
      port map(D => \U1/N_1790\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[25]\);
    
    \U1/cnt_63_0\ : NOR2B
      port map(A => \U1/cnt[0]_net_1\, B => \U1/cnt[1]_net_1\, Y
         => \U1/cnt_63_0_net_1\);
    
    \U1/data_all_RNO_0[105]\ : AO1C
      port map(A => \data_all[105]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[105]\);
    
    \U5/data_send_RNO_23[0]\ : MX2
      port map(A => \data_all[144]\, B => \data_all[152]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_411\);
    
    \U3/data_recive_RNO_1[3]\ : NOR3C
      port map(A => \U3/m36_4\, B => \U3/m36_3\, C => \U3/N_30_0\, 
        Y => \U3/data_recive26\);
    
    \U1/pr_state[6]\ : DFN1C0
      port map(D => \U1/N_256\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U1/pr_state[6]_net_1\);
    
    \U1/data_all_RNO_0[199]\ : AO1C
      port map(A => \data_all[199]\, B => \U1/N_839_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m124_0_i_0\);
    
    \U3/recive_RNO\ : AO1B
      port map(A => \U3/rx_down_net_1\, B => \U3/idle_recive_i_0\, 
        C => \U3/un1_cnt\, Y => \U3/un2_cnt\);
    
    \U1/data_all_RNO_0[196]\ : AO1C
      port map(A => \data_all[196]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m133_i_0_0\);
    
    \U1/data_all_RNO[151]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/m95_1_i_0_0\, Y => \U1/N_130\);
    
    \U5/data_send_RNO_2[0]\ : MX2
      port map(A => \U5/N_459\, B => \U5/N_467\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_515\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I76_Y_0\ : AO1
      port map(A => \U1/N229\, B => \U1/N232\, C => \U1/N227\, Y
         => \U1/ADD_14x14_fast_I76_Y_0\);
    
    \U1/data_all_RNO_0[227]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[227]\, Y => 
        \U1/N_2159\);
    
    \U1/data_all_RNO_0[192]\ : AO1C
      port map(A => \data_all[192]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m145_i_0_0\);
    
    \U1/data_all[234]\ : DFN1E0C0
      port map(D => \U1/N_304\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[234]\);
    
    \U0/sts_ris2\ : DFN1C0
      port map(D => \U0/sts_ris1_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U0/sts_ris2_net_1\);
    
    \U1/data_all_RNO_1[87]\ : NOR2
      port map(A => \U1/data_filter[7]_net_1\, B => \U1/N_834_0\, 
        Y => \U1/N_2136\);
    
    \U1/data_all_RNO_0[23]\ : AO1C
      port map(A => \data_all[23]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m144_0_i_0_0\);
    
    \U1/data_all_RNO[92]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1035\, C
         => \U1/N_1036\, Y => \U1/N_199\);
    
    \U5/data_send_RNO_16[4]\ : MX2
      port map(A => \data_all[36]\, B => \data_all[44]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_359\);
    
    \U0/pr_state_RNI2GH[3]\ : OR2
      port map(A => \U0/pr_state[3]_net_1\, B => 
        \U0/pr_state[5]_net_1\, Y => \U0/N_144\);
    
    \U3/cnt_RNIEAUG_0[2]\ : NOR2
      port map(A => \U3/cnt[2]_net_1\, B => \U3/cnt[6]_net_1\, Y
         => \U3/m41_0\);
    
    \U1/data_all_RNO_0[198]\ : AO1C
      port map(A => \data_all[198]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m127_i_0_0\);
    
    \U5/data_send_RNO_25[6]\ : MX2
      port map(A => \data_all[182]\, B => \data_all[190]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_433\);
    
    \U5/data_send_RNO_20[0]\ : MX2
      port map(A => \data_all[96]\, B => \data_all[104]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_387\);
    
    \U1/data_all_RNO_0[233]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[233]\, Y => 
        \U1/N_911\);
    
    \U1/data_all_RNO[26]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/m135_0_i_0_0\, Y => \U1/N_1791\);
    
    \U1/data_all_RNO[105]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[105]\, Y => \U1/N_1612\);
    
    \U5/data_send_RNO_25[3]\ : MX2
      port map(A => \data_all[179]\, B => \data_all[187]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_430\);
    
    \U1/data_all[61]\ : DFN1E0C0
      port map(D => \U1/N_356\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[61]\);
    
    \U2/parity_check_RNO_7\ : XOR2
      port map(A => \data_send[7]\, B => \U2/parity_check_net_1\, 
        Y => \U2/N_60_i\);
    
    \U2/cnt_RNISS7J_1[1]\ : NOR2B
      port map(A => \U2/N_128\, B => \U2/N_125\, Y => \U2/N_181\);
    
    \U1/data_all[67]\ : DFN1E0C0
      port map(D => \U1/N_169\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[67]\);
    
    \U1/pr_state_0[5]\ : DFN1C0
      port map(D => \U1/N_119\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U1/pr_state_0[5]_net_1\);
    
    \U1/data_all_RNO_0[130]\ : AO1C
      port map(A => \data_all[130]\, B => \U1/N_841_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m205_0_i_0\);
    
    \U5/data_send_RNO_19[1]\ : MX2
      port map(A => \data_all[81]\, B => \data_all[89]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_380\);
    
    \U5/vld_send\ : DFN1E0C0
      port map(D => \U5/pr_state[0]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/N_78\, Q => vld_send);
    
    \rx_uart_pad/U0/U0\ : IOPAD_IN
      port map(PAD => rx_uart, Y => \rx_uart_pad/U0/NET1\);
    
    \U2/cnt_RNI7DUF2_2[10]\ : NOR2B
      port map(A => \U2/N_197\, B => \U2/N_168\, Y => 
        \U2/parity_check_6_sqmuxa\);
    
    \U5/data_send_RNO_16[6]\ : MX2
      port map(A => \data_all[38]\, B => \data_all[46]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_361\);
    
    \U1/data_all_RNO_0[231]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[231]\, Y => 
        \U1/N_985\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I77_Y\ : AO1
      port map(A => \U1/ADD_14x14_fast_I77_un1_Y_0\, B => 
        \U1/N273\, C => \U1/ADD_14x14_fast_I77_Y_2\, Y => 
        \U1/N315\);
    
    \U1/data_all_RNO_0[109]\ : AO1C
      port map(A => \data_all[109]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[109]\);
    
    \U1/cnt_daly_RNO_0[12]\ : OR2B
      port map(A => \U1/m20_N_13_mux\, B => 
        \U1/cnt_daly[11]_net_1\, Y => \U1/N_859\);
    
    \U0/data_ad[2]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[2]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[2]\);
    
    \U2/cnt_n4\ : NOR2B
      port map(A => \U2/cnt_0_sqmuxa_net_1\, B => 
        \U2/cnt_n4_tz_net_1\, Y => \U2/cnt_n4_net_1\);
    
    \U1/data_all_RNO_0[106]\ : AO1C
      port map(A => \data_all[106]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[106]\);
    
    \U5/data_send_RNO_6[6]\ : MX2
      port map(A => \U5/N_345\, B => \U5/N_353\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_465\);
    
    \U4/nx_state[0]\ : DLN0P1C1
      port map(D => \GND\, G => \U4/N_24\, PRE => 
        \U4/nx_state_RNO_0[0]_net_1\, CLR => 
        \U4/nx_state_RNO[0]_net_1\, Q => \U4/nx_state[0]_net_1\);
    
    \U1/data_all_RNO_0[171]\ : AO1C
      port map(A => \data_all[171]\, B => \U1/N_838_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m161_i_0_0\);
    
    \U1/cnt_n2\ : XA1B
      port map(A => \U1/cnt_63_0_net_1\, B => \U1/cnt[2]_net_1\, 
        C => \U1/pr_state_0[7]_net_1\, Y => \U1/cnt_n2_net_1\);
    
    \U1/data_all_RNO_0[102]\ : AO1C
      port map(A => \data_all[102]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[102]\);
    
    \U1/data_all_RNO[229]\ : OA1B
      port map(A => \U1/N_837_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m89_i_0_0\, Y => \U1/N_217\);
    
    \U1/data_all[224]\ : DFN1E0C0
      port map(D => \U1/N_34\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[224]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I44_Y\ : AO1
      port map(A => \U1/N240\, B => \U1/N237\, C => \U1/N236\, Y
         => \U1/N263\);
    
    \U0/rc\ : DFN1E0P0
      port map(D => \U0/N_144\, CLK => sys_clk_c, PRE => 
        sys_rest_c, E => \U0/N_136\, Q => rc_c);
    
    \U1/data_all_RNO_0[64]\ : AO1C
      port map(A => \data_all[64]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m252_i_0_0\);
    
    \U1/data_all_RNO[13]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[13]\, Y => \U1/N_787\);
    
    \U1/data_all_3_0_a2_i_0_o2_0[239]\ : OR3C
      port map(A => \addr_c_0[0]\, B => \U1/I_5_0\, C => 
        \U1/I_9_0\, Y => \U1/m146_i_0_o2_1\);
    
    \U1/data_all[48]\ : DFN1E0C0
      port map(D => \U1/N_702\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[48]\);
    
    \U1/data_all[156]\ : DFN1E0C0
      port map(D => \U1/N_744\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[156]\);
    
    \U5/data_send_RNO_24[2]\ : MX2
      port map(A => \data_all[162]\, B => \data_all[170]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_421\);
    
    \U5/data_send_RNO_21[1]\ : MX2
      port map(A => \data_all[113]\, B => \data_all[121]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_396\);
    
    \U3/cnt_RNIJFUG[6]\ : NOR2A
      port map(A => \U3/cnt[6]_net_1\, B => \U3/cnt[7]_net_1\, Y
         => \U3/m11_2\);
    
    \U1/cnt_daly_RNIO51Q[12]\ : NOR2A
      port map(A => \U1/cnt_daly[12]_net_1\, B => 
        \U1/cnt_daly[10]_net_1\, Y => \U1/m61_0_i_a3_1_0\);
    
    \U1/data_all_RNO_0[141]\ : AO1C
      port map(A => \data_all[141]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[141]\);
    
    \U1/data_all_RNO_0[108]\ : AO1C
      port map(A => \data_all[108]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[108]\);
    
    \U1/data_all_RNO_0[38]\ : AO1C
      port map(A => \data_all[38]\, B => \U1/N_832\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m280_i_0_0\);
    
    \data_in_pad[2]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[2]/U0/NET1\, Y => 
        \data_in_c[2]\);
    
    \U5/data_send_RNO_23[7]\ : MX2
      port map(A => \data_all[151]\, B => \data_all[159]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_418\);
    
    \U4/conver_ris3\ : DFN1P0
      port map(D => \U4/conver_ris2_i\, CLK => sys_clk_c, PRE => 
        sys_rest_c, Q => \U4/conver_ris3_i_0\);
    
    \U5/data_send_RNO_14[7]\ : MX2
      port map(A => \data_all[7]\, B => \data_all[15]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_346\);
    
    \U1/data_all_3_i_0_0_o2_1[190]\ : OR3B
      port map(A => \U1/I_5_0\, B => \U1/I_9_0\, C => 
        \addr_c_0[0]\, Y => \U1/data_all_3_i_0_0_o2_1[190]_net_1\);
    
    \U1/data_all_RNO_0[24]\ : AO1C
      port map(A => \data_all[24]\, B => \U1/N_836\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m141_0_i_0_0\);
    
    \U1/pr_state_RNO[6]\ : AO1A
      port map(A => \U1/N_860\, B => \U1/N_856\, C => 
        \U1/m77_i_0_0\, Y => \U1/N_256\);
    
    \U1/data_all[143]\ : DFN1E0C0
      port map(D => \U1/N_17\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[143]\);
    
    \U0/data_ad_RNO[5]\ : NOR2A
      port map(A => \data_in_c[5]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[5]\);
    
    \U1/data_all_RNO[124]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[124]\, Y => \U1/N_388\);
    
    \U1/data_all_RNO[221]\ : OA1B
      port map(A => \U1/N_840\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m57_0_i_0_0\, Y => \U1/N_1780\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I8_P0N\ : OR2
      port map(A => \data_ad[8]\, B => \U1/data_filter[8]_net_1\, 
        Y => \U1/N201\);
    
    \U2/cnt_RNIDTJ9[2]\ : NOR2A
      port map(A => \U2/cnt[7]_net_1\, B => \U2/cnt[2]_net_1\, Y
         => \U2/N_124\);
    
    \U1/data_all[163]\ : DFN1E0C0
      port map(D => \U1/N_1816\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[163]\);
    
    \U1/data_filter[11]\ : DFN1E0C0
      port map(D => \U1/N_35\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[11]_net_1\);
    
    \U1/cnt_daly_RNO[10]\ : XA1B
      port map(A => \U1/m22_N_11_mux\, B => 
        \U1/cnt_daly[10]_net_1\, C => \U1/pr_state_0[7]_net_1\, Y
         => \U1/cnt_daly_n10\);
    
    \U1/data_filter[9]\ : DFN1E0C0
      port map(D => \U1/N_46_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[9]_net_1\);
    
    \U2/parity_check_RNO_2\ : AO1A
      port map(A => \U2/N_60_i\, B => \U2/parity_check_8_sqmuxa\, 
        C => \U2/N_116\, Y => \U2/parity_check_10_iv_0_2\);
    
    \U1/data_all_RNO[220]\ : OA1B
      port map(A => \U1/N_840\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[220]\, Y => \U1/N_166\);
    
    \U1/data_all_RNO_0[98]\ : AO1C
      port map(A => \data_all[98]\, B => \U1/N_829_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[98]\);
    
    \U1/data_all_RNO[39]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2205\, C
         => \U1/N_2206\, Y => \U1/N_1812\);
    
    \U1/data_all[42]\ : DFN1E0C0
      port map(D => \U1/N_278\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[42]\);
    
    \U3/cnt_4[11]\ : XA1
      port map(A => \U3/N_2\, B => \U3/cnt[11]_net_1\, C => 
        \U3/recive_net_1\, Y => \U3/cnt_4[11]_net_1\);
    
    \U5/data_send_RNO_23[4]\ : MX2
      port map(A => \data_all[148]\, B => \data_all[156]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_415\);
    
    \U1/data_all_RNO_1[92]\ : NOR2
      port map(A => \U1/data_filter[12]_net_1\, B => \U1/N_834\, 
        Y => \U1/N_1036\);
    
    \U5/cnt_RNI5FPF[0]\ : CLKINT
      port map(A => \U5/cnt_0[0]\, Y => \U5/cnt[0]_net_1\);
    
    \U5/data_send_RNO_2[5]\ : MX2
      port map(A => \U5/N_464\, B => \U5/N_472\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_520\);
    
    \U5/data_send_RNO_23[3]\ : MX2
      port map(A => \data_all[147]\, B => \data_all[155]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_414\);
    
    \U1/data_all_RNO[107]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[11]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[107]\, Y => \U1/N_44\);
    
    \U2/tx_uart_RNO_7\ : AO1
      port map(A => \U2/tx_uart36\, B => \U2/parity_check_net_1\, 
        C => \U2/tx_uart_11_iv_0\, Y => \U2/tx_uart_11_iv_1\);
    
    \U1/data_all_RNO[9]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1077\, C
         => \U1/N_1078\, Y => \U1/N_243\);
    
    \U1/cnt_n0\ : NOR2
      port map(A => \U1/cnt[0]_net_1\, B => 
        \U1/pr_state[7]_net_1\, Y => \U1/N_1415\);
    
    \U1/data_all_RNO[47]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_832\, C
         => \data_all[47]\, Y => \U1/data_all_3[47]\);
    
    \U1/data_filter_RNO_0[1]\ : AO1D
      port map(A => \U1/data_filter[3]_net_1\, B => 
        \U1/pr_state[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, Y
         => \U1/m57_0_0_0\);
    
    \U1/data_all_RNO_0[232]\ : AO1C
      port map(A => \data_all[232]\, B => \U1/N_837_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m82_0_i_0_0\);
    
    \U1/data_all_RNO_0[91]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[91]\, Y => 
        \U1/N_2131\);
    
    \U1/data_all_RNO[119]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[119]\, Y => \U1/N_378\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I30_Y\ : AO1
      port map(A => \U1/N182\, B => \U1/N186\, C => \U1/N185\, Y
         => \U1/N246\);
    
    \U1/data_all_RNO_0[209]\ : NOR2A
      port map(A => \U1/N_840\, B => \data_all[209]\, Y => 
        \U1/N_1031\);
    
    \U1/data_all_RNO_0[163]\ : AO1C
      port map(A => \data_all[163]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m185_i_0_0\);
    
    \U1/data_all_RNO[95]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_834_0\, C
         => \data_all[95]\, Y => \U1/data_all_3[95]\);
    
    \U0/pr_state[3]\ : DFN1C0
      port map(D => \U0/pr_state_ns[2]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U0/pr_state[3]_net_1\);
    
    \U1/data_all[159]\ : DFN1E0C0
      port map(D => \U1/data_all_3[159]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[159]\);
    
    \U1/data_all[187]\ : DFN1E0C0
      port map(D => \U1/N_415\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[187]\);
    
    \U1/data_all_RNO_0[220]\ : AO1C
      port map(A => \data_all[220]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[220]\);
    
    \U1/data_all_RNO_0[154]\ : AO1C
      port map(A => \data_all[154]\, B => \U1/N_842_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m88_0_i_0_0\);
    
    \U2/cnt_RNIOOHD2[5]\ : NOR2B
      port map(A => \U2/tx_uart38_1\, B => \U2/tx_uart38_10\, Y
         => \U2/tx_uart38\);
    
    \U1/delay_channel1_RNO\ : AO1
      port map(A => \U1/m101_i_0_a3_0_0\, B => \U4.N_31\, C => 
        \U1/N_872\, Y => \U1/N_1838\);
    
    \data_in_pad[6]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[6]/U0/NET1\, Y => 
        \data_in_c[6]\);
    
    \U5/data_send_RNO_23[5]\ : MX2
      port map(A => \data_all[149]\, B => \data_all[157]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_416\);
    
    \U1/data_all[29]\ : DFN1E0C0
      port map(D => \U1/N_763\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[29]\);
    
    \U2/cnt_n6\ : NOR2B
      port map(A => \U2/cnt_0_sqmuxa_net_1\, B => 
        \U2/cnt_n6_tz_net_1\, Y => \U2/cnt_n6_net_1\);
    
    \U1/data_all_RNO_0[48]\ : AO1C
      port map(A => \data_all[48]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[48]\);
    
    \U1/data_all_RNO_0[167]\ : AO1C
      port map(A => \data_all[167]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m173_i_0_0\);
    
    \U5/data_send_RNO_18[6]\ : MX2
      port map(A => \data_all[70]\, B => \data_all[78]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_377\);
    
    \U4/conver_ris_RNIE5931\ : NOR3B
      port map(A => \U4.N_31\, B => \U4/conver_ris_net_1\, C => 
        \addr_c_0[0]\, Y => \U4/N_22\);
    
    \U2/cnt_RNINV8G1[3]\ : NOR3C
      port map(A => \U2/tx_uart37_1\, B => \U2/tx_uart37_0\, C
         => \U2/tx_uart37_6_0\, Y => \U2/tx_uart37_8\);
    
    \U2/cnt_RNI9QRS[1]\ : NOR3C
      port map(A => \U2/N_125\, B => \U2/N_124\, C => \U2/N_163\, 
        Y => \U2/N_196\);
    
    \U1/data_all_RNO[12]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[12]\, Y => \U1/N_239\);
    
    \U1/cnt_daly_RNO_1[9]\ : NOR3C
      port map(A => \U1/cnt_daly[4]_net_1\, B => 
        \U1/cnt_daly[6]_net_1\, C => \U1/m24_m4_e_2\, Y => 
        \U1/m24_m4_e_4\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I71_un1_Y\ : NOR3C
      port map(A => \U1/N245\, B => \U1/N249\, C => \U1/N176\, Y
         => \U1/I71_un1_Y\);
    
    \U5/data_send_RNO_0[6]\ : MX2C
      port map(A => \U5/N_521\, B => \U5/N_529\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i71_mux\);
    
    \U1/data_all_RNO_0[77]\ : AO1C
      port map(A => \data_all[77]\, B => \U1/N_833\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m212_0_i_0\);
    
    \U0/cnt_rc_n1\ : XA1B
      port map(A => \U0/cnt_rc[1]_net_1\, B => 
        \U0/cnt_rc[0]_net_1\, C => \U0/pr_state[4]_net_1\, Y => 
        \U0/cnt_rc_n1_net_1\);
    
    \U3/cnt_RNIJIC91[1]\ : NOR3B
      port map(A => \U3/cnt[0]_net_1\, B => \U3/m11_4\, C => 
        \U3/cnt[1]_net_1\, Y => \U3/m11_8\);
    
    \U1/data_all_RNO[41]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/m271_i_0_0\, Y => \U1/N_272\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I29_Y\ : NOR2B
      port map(A => \U1/N186\, B => \U1/N189\, Y => \U1/N245\);
    
    \U1/m107_e\ : NOR3C
      port map(A => \U1/m107_e_2_net_1\, B => \U1/m107_e_1_net_1\, 
        C => \U1/m107_e_3_net_1\, Y => \U1/N_139\);
    
    \U1/data_all[41]\ : DFN1E0C0
      port map(D => \U1/N_272\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[41]\);
    
    \U5/data_send_RNO_5[1]\ : MX2
      port map(A => \U5/N_508\, B => \U5/N_67_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_68\);
    
    \U5/data_send_RNO_15[1]\ : MX2
      port map(A => \data_all[17]\, B => \data_all[25]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_348\);
    
    \U1/data_all_RNO_0[41]\ : AO1C
      port map(A => \data_all[41]\, B => \U1/N_832\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m271_i_0_0\);
    
    \U1/data_filter_RNO[12]\ : XA1
      port map(A => \U1/data_filter[12]_net_1\, B => \U1/N315\, C
         => \U1/pr_state_0[5]_net_1\, Y => \U1/data_filter_4[12]\);
    
    \U1/data_all_RNO_1[75]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_833\, 
        Y => \U1/N_958\);
    
    \U1/data_all[47]\ : DFN1E0C0
      port map(D => \U1/data_all_3[47]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[47]\);
    
    \U1/data_all_RNO[57]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2143\, C
         => \U1/N_2144\, Y => \U1/N_688\);
    
    \U1/data_all_RNO[149]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m103_0_i_0_0\, Y => \U1/N_1797\);
    
    \U5/data_send_RNO_6[2]\ : MX2
      port map(A => \U5/N_341\, B => \U5/N_349\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_461\);
    
    \U5/data_send_RNO_12[2]\ : MX2
      port map(A => \U5/N_437\, B => \U5/N_445\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_509\);
    
    \U2/cnt_RNIOO7J[1]\ : NOR3C
      port map(A => \U2/cnt[7]_net_1\, B => \U2/cnt[1]_net_1\, C
         => \U2/un1_cnt_4\, Y => \U2/tx_uart34_0_a2_2_2\);
    
    \U1/data_all_RNO[74]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_959\, C
         => \U1/N_960\, Y => \U1/N_183\);
    
    \U1/cnt[1]\ : DFN1E1C0
      port map(D => \U1/cnt_n1_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_793\, Q => \U1/cnt[1]_net_1\);
    
    \U1/data_all_RNO_0[2]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[2]\, Y => 
        \U1/N_981\);
    
    \U5/data_send_RNO_6[4]\ : MX2
      port map(A => \U5/N_343\, B => \U5/N_351\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_463\);
    
    \U4/nx_state_RNO_0[0]\ : MX2
      port map(A => \U4/N_27\, B => \U4/N_25\, S => 
        \U4/pr_state[0]_net_1\, Y => \U4/nx_state_RNO_0[0]_net_1\);
    
    \U0/sts_ris1\ : DFN1C0
      port map(D => sts_c, CLK => sys_clk_c, CLR => sys_rest_c, Q
         => \U0/sts_ris1_net_1\);
    
    \U5/data_send_RNO_7[4]\ : MX2
      port map(A => \U5/N_359\, B => \U5/N_367\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_471\);
    
    \U3/un7_cnt_1_I_22\ : AND3
      port map(A => \U3/DWACT_FINC_E[0]\, B => 
        \U3/DWACT_FINC_E[2]\, C => \U3/DWACT_FINC_E[3]\, Y => 
        \U3/N_5\);
    
    \U3/un7_cnt_1_I_12\ : AX1C
      port map(A => \U3/cnt[3]_net_1\, B => \U3/DWACT_FINC_E[0]\, 
        C => \U3/cnt[4]_net_1\, Y => \U3/I_12\);
    
    \U1/data_all[197]\ : DFN1E0C0
      port map(D => \U1/N_89\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[197]\);
    
    \U5/data_send_RNO_9[0]\ : MX2
      port map(A => \U5/N_387\, B => \U5/N_395\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_483\);
    
    \U1/data_all_RNO_1[39]\ : NOR2
      port map(A => \U1/data_filter[7]_net_1\, B => \U1/N_832\, Y
         => \U1/N_2206\);
    
    \U5/cnt_RNIBVIV[1]\ : NOR2B
      port map(A => \U5/cnt[1]_net_1\, B => \U5/cnt[0]_net_1\, Y
         => \U5/N_10_0\);
    
    \U2/cnt_n3\ : XA1
      port map(A => \U2/cnt_c2_net_1\, B => \U2/cnt[3]_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n3_net_1\);
    
    \addr_pad[3]/U0/U0\ : IOPAD_TRI
      port map(D => \addr_pad[3]/U0/NET1\, E => 
        \addr_pad[3]/U0/NET2\, PAD => addr(3));
    
    \U5/data_send_RNO_21[7]\ : MX2
      port map(A => \data_all[119]\, B => \data_all[127]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_402\);
    
    \U5/data_send_RNO_20[4]\ : MX2
      port map(A => \data_all[100]\, B => \data_all[108]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_391\);
    
    \ce_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => ce_c, E => \VCC\, DOUT => \ce_pad/U0/NET1\, 
        EOUT => \ce_pad/U0/NET2\);
    
    \U3/idle_recive\ : DFN1P0
      port map(D => \U3/recive_i\, CLK => sys_clk_c, PRE => 
        sys_rest_c, Q => \U3/idle_recive_i_0\);
    
    \U3/data_recive_RNO[4]\ : MX2
      port map(A => \U3/m85_0\, B => rx_uart_c, S => 
        \U3/data_recive27\, Y => \U3/data_recive_12[4]\);
    
    \U5/data_send_RNO_1[4]\ : MX2A
      port map(A => \U5/N_533\, B => \U5/N_47_0\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_48_0\);
    
    \U2/cnt_c1_i_RNI3JEJ\ : AND3B
      port map(A => \U2/cnt[2]_net_1\, B => \U2/N_7\, C => 
        \U2/cnt[8]_net_1\, Y => \U2/tx_uart38_10_4\);
    
    \U1/data_all[116]\ : DFN1E0C0
      port map(D => \U1/N_372\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[116]\);
    
    \U2/cnt_RNIH1K9_0[9]\ : NOR2A
      port map(A => \U2/cnt[9]_net_1\, B => \U2/cnt[4]_net_1\, Y
         => \U2/N_164\);
    
    \U5/cnt[1]\ : DFN1E0C0
      port map(D => \U5/cnt_n1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \U5/cnt_0[1]\);
    
    \U3/cnt_RNIMLC91[2]\ : NOR2A
      port map(A => \U3/N_29\, B => \U3/cnt[2]_net_1\, Y => 
        \U3/N_30_0\);
    
    \U1/data_all_RNO[84]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1043\, C
         => \U1/N_1044\, Y => \U1/N_210\);
    
    \U2/cnt_n9\ : XA1
      port map(A => \U2/cnt_c8_net_1\, B => \U2/cnt[9]_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n9_net_1\);
    
    \U5/data_send_RNO_18[0]\ : MX2
      port map(A => \data_all[64]\, B => \data_all[72]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_371\);
    
    \U4/addr_0[0]\ : DFN1E0C0
      port map(D => \U4/N_20\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U4/N_7_0\, Q => \addr_c_0[0]\);
    
    \U1/data_all_RNO_0[203]\ : AO1C
      port map(A => \data_all[203]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m112_0_0_i_0\);
    
    \U1/data_all_RNO[51]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2151\, C
         => \U1/N_2152\, Y => \U1/N_696\);
    
    \data_in_pad[8]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(8), Y => \data_in_pad[8]/U0/NET1\);
    
    \U5/data_send_RNO_15[5]\ : MX2
      port map(A => \data_all[21]\, B => \data_all[29]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_352\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I2_P0N\ : OR2
      port map(A => \data_ad[2]\, B => \U1/data_filter[2]_net_1\, 
        Y => \U1/N183\);
    
    \U5/data_send_RNO_6[1]\ : MX2
      port map(A => \U5/N_340\, B => \U5/N_348\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_460\);
    
    \U1/data_all_RNO_0[75]\ : NOR2A
      port map(A => \U1/N_833\, B => \data_all[75]\, Y => 
        \U1/N_957\);
    
    \U0/data_ad[4]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[4]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[4]\);
    
    \U1/data_all_RNO_1[1]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_835\, Y
         => \U1/N_1099\);
    
    \U1/data_all_RNO[166]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/m176_i_0_0\, Y => \U1/N_319\);
    
    \U1/m253_i_0_o2_0\ : OR3B
      port map(A => \U1/I_5_0\, B => \addr_c[0]\, C => \U1/I_9_0\, 
        Y => \U1/m253_i_0_o2_0_net_1\);
    
    \U5/data_send_RNO_4[0]\ : MX2C
      port map(A => \U5/N_491\, B => \U5/N_499\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_537\);
    
    \U1/data_all_RNO_1[211]\ : NOR2
      port map(A => \U1/data_filter[3]_net_1\, B => \U1/N_840\, Y
         => \U1/N_1030\);
    
    \U1/data_all[140]\ : DFN1E0C0
      port map(D => \U1/N_94\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[140]\);
    
    \U1/data_all_RNO_0[100]\ : AO1C
      port map(A => \data_all[100]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[100]\);
    
    \U1/data_all[84]\ : DFN1E0C0
      port map(D => \U1/N_210\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[84]\);
    
    \U5/data_send_RNO_16[5]\ : MX2
      port map(A => \data_all[37]\, B => \data_all[45]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_360\);
    
    \U5/cnt_RNO[0]\ : NOR2A
      port map(A => \U5/pr_state[1]_net_1\, B => 
        \U5/cnt[0]_net_1\, Y => \U5/N_21_0\);
    
    \U2/cnt_RNIH1K9[9]\ : NOR2A
      port map(A => \U2/cnt[4]_net_1\, B => \U2/cnt[9]_net_1\, Y
         => \U2/N_125\);
    
    \U1/data_all_RNO[36]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/m286_i_0_0\, Y => \U1/N_1809\);
    
    \U1/data_all[160]\ : DFN1E0C0
      port map(D => \U1/N_1814\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[160]\);
    
    \U1/data_all_RNO_0[201]\ : AO1C
      port map(A => \data_all[201]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m118_0_i_0_0\);
    
    \U5/data_send_RNO_20[2]\ : MX2
      port map(A => \data_all[98]\, B => \data_all[106]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_389\);
    
    \U1/data_all_RNO_0[125]\ : AO1C
      port map(A => \data_all[125]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[125]\);
    
    \U1/m146_i_0_o2_0\ : OR2
      port map(A => \U1/I_7_0\, B => \U1/OVER\, Y => \U1/N_817\);
    
    \U1/data_all[80]\ : DFN1E0C0
      port map(D => \U1/N_224\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[80]\);
    
    \U1/data_filter[7]\ : DFN1E0C0
      port map(D => \U1/N_49_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[7]_net_1\);
    
    \U5/data_send_RNO_4[2]\ : MX2C
      port map(A => \U5/N_493\, B => \U5/N_501\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_535\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I49_Y\ : NOR2B
      port map(A => \U1/N241\, B => \U1/N245\, Y => \U1/N268\);
    
    \U2/cnt_RNIK3R61[9]\ : NOR3C
      port map(A => \U2/cnt[0]_net_1\, B => \U2/cnt[9]_net_1\, C
         => \U2/N_177\, Y => \U2/tx_uart36_6\);
    
    \U3/cnt[9]\ : DFN1C0
      port map(D => \U3/I_26\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/cnt[9]_net_1\);
    
    \U0/cnt_rc[3]\ : DFN1E0C0
      port map(D => \U0/cnt_rc_n3_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U0/N_135\, Q => 
        \U0/cnt_rc[3]_net_1\);
    
    \U2/cnt_RNIETQ61_0[0]\ : NOR2B
      port map(A => \U2/N_177\, B => \U2/N_126\, Y => 
        \U2/tx_uart34_1\);
    
    \U1/data_all_RNO[64]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/m252_i_0_0\, Y => \U1/N_163\);
    
    \U2/cnt_RNIBRJ9_0[1]\ : NOR2A
      port map(A => \U2/cnt[6]_net_1\, B => \U2/cnt[1]_net_1\, Y
         => \U2/N_128\);
    
    \U1/data_all_RNO[225]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2163\, C
         => \U1/N_2164\, Y => \U1/N_708\);
    
    \U1/data_all[219]\ : DFN1E0C0
      port map(D => \U1/N_170\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[219]\);
    
    \U1/data_all[175]\ : DFN1E0C0
      port map(D => \U1/data_all_3[175]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[175]\);
    
    \sys_rest_pad/U0/U1\ : CLKIO
      port map(A => \sys_rest_pad/U0/NET1\, Y => sys_rest_c);
    
    \U1/data_all[86]\ : DFN1E0C0
      port map(D => \U1/N_205\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[86]\);
    
    \U2/tx_uart_RNO_2\ : AO1
      port map(A => \U2/parity_check_1_sqmuxa\, B => 
        \data_send[0]\, C => \U2/data_send_m[2]\, Y => 
        \U2/tx_uart_11_iv_5\);
    
    \U1/data_all_RNO_0[134]\ : AO1C
      port map(A => \data_all[134]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[134]\);
    
    \U1/data_all_RNO[176]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[176]\, Y => \U1/N_393\);
    
    \U2/parity_check_RNO_16\ : XOR2
      port map(A => \data_send[3]\, B => \U2/parity_check_net_1\, 
        Y => \U2/N_59_i\);
    
    \U5/data_send_RNO_7[0]\ : MX2
      port map(A => \U5/N_355\, B => \U5/N_363\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_467\);
    
    \U1/data_filter_RNO_0[3]\ : AO1D
      port map(A => \U1/data_filter[5]_net_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, 
        Y => \U1/data_filter_4_i_0_0_0[3]\);
    
    \U1/data_all[106]\ : DFN1E0C0
      port map(D => \U1/N_46\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[106]\);
    
    \U2/cnt_RNI8O7O[9]\ : NOR3A
      port map(A => \U2/cnt[11]_net_1\, B => \U2/cnt[9]_net_1\, C
         => \U2/cnt[7]_net_1\, Y => \U2/un1_cnt_5\);
    
    \U1/data_all_RNO[128]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[128]\, Y => \U1/N_1835\);
    
    \U5/data_send_RNO_14[0]\ : MX2
      port map(A => \data_all[0]\, B => \data_all[8]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_339\);
    
    \U2/cnt_RNITKMOB[10]\ : OR3
      port map(A => \U2/un1_tx_uart27_4\, B => 
        \U2/un1_tx_uart27_0\, C => \U2/un1_tx_uart27_4_1\, Y => 
        \U2/un1_tx_uart27_5\);
    
    \U1/data_all_RNO[15]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_835_0\, C
         => \data_all[15]\, Y => \U1/data_all_3[15]\);
    
    \U1/data_all[119]\ : DFN1E0C0
      port map(D => \U1/N_378\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[119]\);
    
    \U1/data_all_RNO[163]\ : OA1B
      port map(A => \U1/N_838\, B => \U1/data_filter[3]_net_1\, C
         => \U1/m185_i_0_0\, Y => \U1/N_1816\);
    
    \U0/data_ad_RNO[6]\ : NOR2A
      port map(A => \data_in_c[6]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[6]\);
    
    \U1/data_all_RNO[156]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/m82_1_i_i_0\, Y => \U1/N_744\);
    
    \U1/data_all_RNO[160]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/m191_i_0_0\, Y => \U1/N_1814\);
    
    \U1/data_all_RNO[209]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1031\, C
         => \U1/N_1032\, Y => \U1/N_194\);
    
    \U1/data_all[85]\ : DFN1E0C0
      port map(D => \U1/N_208\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[85]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I71_Y\ : OR2
      port map(A => \U1/I71_un1_Y\, B => \U1/N271\, Y => 
        \U1/N332\);
    
    \U5/data_send_RNO_4[7]\ : MX2C
      port map(A => \U5/N_498\, B => \U5/N_506\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_530\);
    
    \U5/cnt[0]\ : DFN1E0C0
      port map(D => \U5/N_21_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \U5/cnt_0[0]\);
    
    \U1/data_filter_RNO[4]\ : OA1C
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/un2_data_filter[4]\, C => 
        \U1/data_filter_4_i_0_0_0[4]\, Y => \U1/N_41\);
    
    \U1/data_all_RNO_0[129]\ : AO1C
      port map(A => \data_all[129]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[129]\);
    
    \U2/cnt_RNIQRF61[1]\ : NOR3C
      port map(A => \U2/N_176\, B => \U2/N_129\, C => 
        \U2/tx_uart34_0_a2_2_2\, Y => \U2/N_194\);
    
    \U1/data_all[14]\ : DFN1E0C0
      port map(D => \U1/data_all_3[14]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[14]\);
    
    \U5/data_send_RNO_11[3]\ : MX2
      port map(A => \U5/N_422\, B => \U5/N_430\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_502\);
    
    \U1/pr_state_RNO_1[3]\ : NOR3A
      port map(A => ad_over, B => \U1/pr_state[3]_net_1\, C => 
        \U1/N_854\, Y => \U1/N_870\);
    
    \U1/pr_state_RNINLAR[6]\ : NOR2B
      port map(A => ad_over, B => \U1/pr_state[6]_net_1\, Y => 
        \U1/N_119\);
    
    \U1/cnt_daly[0]\ : DFN1E0C0
      port map(D => \U1/N_42\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[0]_net_1\);
    
    \U1/m79_0_i_i_o2_0_0\ : OR2
      port map(A => \U1/m79_0_i_i_o2_0_net_1\, B => \U1/N_817\, Y
         => \U1/N_842_0\);
    
    \U1/data_all_RNO_0[122]\ : AO1C
      port map(A => \data_all[122]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[122]\);
    
    \U1/cnt_daly_RNISPUL1[4]\ : NOR3A
      port map(A => \U1/m24_m4_e_2\, B => \U1/cnt_daly[5]_net_1\, 
        C => \U1/cnt_daly[4]_net_1\, Y => \U1/m61_0_i_a3_1_8\);
    
    \U1/receive_on_RNO_0\ : NOR3B
      port map(A => \U1/cnt_receive_over_net_1\, B => 
        \U1/receive_flag_net_1\, C => \data_recive[0]\, Y => 
        \U1/m110_i_0_a3_1\);
    
    \U1/data_all_RNO[104]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[104]\, Y => \U1/N_50\);
    
    \U5/data_send_RNO_5[7]\ : MX2
      port map(A => \U5/N_514\, B => \U5/N_25_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_26_0\);
    
    \U5/data_send_RNO_15[2]\ : MX2
      port map(A => \data_all[18]\, B => \data_all[26]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_349\);
    
    \U1/data_all_RNO_0[202]\ : NOR2A
      port map(A => \U1/N_839\, B => \data_all[202]\, Y => 
        \U1/N_925\);
    
    \U1/data_all_RNO[201]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/m118_0_i_0_0\, Y => \U1/N_2041\);
    
    \U1/data_all[10]\ : DFN1E0C0
      port map(D => \U1/N_789\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[10]\);
    
    \U5/data_send_RNO_8[0]\ : MX2
      port map(A => \U5/N_371\, B => \U5/N_379\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_475\);
    
    \U5/cnt_RNO[3]\ : XA1
      port map(A => \U5/cnt[3]_net_1\, B => \U5/N_11_0\, C => 
        \U5/pr_state[1]_net_1\, Y => \U5/cnt_n3\);
    
    \U4/addr_RNIE18V[3]\ : NOR2B
      port map(A => \U4/N_9_0\, B => \addr_c[3]\, Y => 
        \U4/N_10_0\);
    
    \U2/cnt_RNICSJ9[2]\ : NOR2B
      port map(A => \U2/cnt[2]_net_1\, B => \U2/cnt[6]_net_1\, Y
         => \U2/un1_cnt_4\);
    
    \U1/data_all_RNO_0[90]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[90]\, Y => 
        \U1/N_2291\);
    
    \U1/data_all_3_i_0_0_o2[190]\ : OR2
      port map(A => \U1/data_all_3_i_0_0_o2_1[190]_net_1\, B => 
        \U1/N_817\, Y => \U1/N_844\);
    
    \U1/data_all[183]\ : DFN1E0C0
      port map(D => \U1/N_407\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[183]\);
    
    \U0/pr_state_RNO[5]\ : MX2
      port map(A => \U0/pr_state[1]_net_1\, B => 
        \U0/conver_ris_i_0\, S => \U0/pr_state[5]_net_1\, Y => 
        \U0/pr_state_ns[0]\);
    
    \U1/data_all_RNO_0[128]\ : AO1C
      port map(A => \data_all[128]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[128]\);
    
    \U1/data_all_RNO_1[42]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_832\, 
        Y => \U1/N_2200\);
    
    \U4/conver_ris1\ : DFN1C0
      port map(D => receive_on, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U4/conver_ris1_net_1\);
    
    \data_in_pad[3]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[3]/U0/NET1\, Y => 
        \data_in_c[3]\);
    
    \U5/data_send_RNO_12[3]\ : MX2
      port map(A => \U5/N_438\, B => \U5/N_446\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_510\);
    
    \U1/data_all[137]\ : DFN1E0C0
      port map(D => \U1/N_87\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[137]\);
    
    \U1/cnt_daly_RNO[5]\ : XA1C
      port map(A => \U1/cnt_daly[5]_net_1\, B => \U1/N_848\, C
         => \U1/pr_state[7]_net_1\, Y => \U1/N_804\);
    
    \U1/cnt_daly_RNI3K9S5[1]\ : NOR3C
      port map(A => \U1/m61_0_i_a3_1_8\, B => \U1/m61_0_i_a3_1_7\, 
        C => \U1/m61_0_i_a3_1_9\, Y => \U1/N_866\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I94_Y\ : XOR3
      port map(A => \U1/data_filter[6]_net_1\, B => \data_ad[6]\, 
        C => \U1/N329\, Y => \U1/un2_data_filter[6]\);
    
    \U1/data_all_RNO[173]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m153_i_0_0\, Y => \U1/N_333\);
    
    \U1/data_all[54]\ : DFN1E0C0
      port map(D => \U1/N_43\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[54]\);
    
    \U1/data_all[209]\ : DFN1E0C0
      port map(D => \U1/N_194\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[209]\);
    
    \U1/data_all_RNO[170]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/m164_i_0_0\, Y => \U1/N_327\);
    
    \U1/cnt_daly_RNO[11]\ : XA1B
      port map(A => \U1/cnt_daly[11]_net_1\, B => 
        \U1/m20_N_13_mux\, C => \U1/pr_state[7]_net_1\, Y => 
        \U1/cnt_daly_n11\);
    
    \U1/data_all_RNO[200]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/m121_0_0_i_0\, Y => \U1/N_2042\);
    
    \U1/data_all[16]\ : DFN1E0C0
      port map(D => \U1/N_1782\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[16]\);
    
    \U5/data_send_RNO_24[3]\ : MX2
      port map(A => \data_all[163]\, B => \data_all[171]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_422\);
    
    \U3/data_recive_RNO_2[6]\ : NOR3A
      port map(A => \U3/m79_2\, B => \U3/cnt[8]_net_1\, C => 
        \U3/cnt[5]_net_1\, Y => \U3/m79_4\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I55_Y\ : AO1
      port map(A => \U1/N249\, B => \U1/N176\, C => \U1/N248\, Y
         => \U1/N275\);
    
    \U5/cnt_RNO[4]\ : XA1
      port map(A => \U5/cnt[4]_net_1\, B => \U5/N_12_0\, C => 
        \U5/pr_state[1]_net_1\, Y => \U5/cnt_n4\);
    
    \U1/data_all_RNO_0[58]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[58]\, Y => 
        \U1/N_2141\);
    
    \U1/data_all_RNO[153]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2231\, C
         => \U1/N_2232\, Y => \U1/N_1799\);
    
    \U1/data_all[50]\ : DFN1E0C0
      port map(D => \U1/N_698\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[50]\);
    
    \U1/m103_i_o2_0_o2_0\ : OR2
      port map(A => \U1/m103_i_o2_0_o2_0_net_1\, B => \U1/N_818\, 
        Y => \U1/N_839_0\);
    
    \U1/data_all_3_i_0_0_o2[111]\ : OR3A
      port map(A => \addr_c_0[0]\, B => \U1/N_818\, C => 
        \U1/N_820\, Y => \U1/N_829\);
    
    \U1/data_all[109]\ : DFN1E0C0
      port map(D => \U1/N_1610\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[109]\);
    
    \U1/data_all_RNO_0[151]\ : AO1C
      port map(A => \data_all[151]\, B => \U1/N_842_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m95_1_i_0_0\);
    
    \U1/data_all_RNO[150]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/m98_0_i_i_0\, Y => \U1/N_751\);
    
    \U1/data_all_RNO_1[28]\ : NOR2
      port map(A => \U1/data_filter[12]_net_1\, B => \U1/N_836\, 
        Y => \U1/N_2254\);
    
    \U1/cnt[0]\ : DFN1E1C0
      port map(D => \U1/N_1415\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_793\, Q => \U1/cnt[0]_net_1\);
    
    \U1/cnt_daly_RNO[12]\ : XA1C
      port map(A => \U1/cnt_daly[12]_net_1\, B => \U1/N_859\, C
         => \U1/pr_state_0[7]_net_1\, Y => \U1/cnt_daly_n12\);
    
    \U0/cnt_rc_RNI9BJE[3]\ : NOR3B
      port map(A => \U0/pr_state[0]_net_1\, B => 
        \U0/cnt_rc[3]_net_1\, C => \U0/cnt_rc[1]_net_1\, Y => 
        \U0/pr_state_ns_a4_2[1]\);
    
    \U1/data_all_RNO[99]\ : OA1B
      port map(A => \U1/N_829\, B => \U1/data_filter[3]_net_1\, C
         => \U1/data_all_3_i_0_0_0[99]\, Y => \U1/N_60\);
    
    \U1/cnt_daly[9]\ : DFN1E0C0
      port map(D => \U1/cnt_daly_n9\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[9]_net_1\);
    
    \U1/data_all_RNO_0[40]\ : AO1C
      port map(A => \data_all[40]\, B => \U1/N_832\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m274_i_0_0\);
    
    \U2/cnt_24_0\ : NOR2B
      port map(A => \U2/cnt[10]_net_1\, B => 
        \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_24_0_net_1\);
    
    \U1/data_all_RNO[40]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/m274_i_0_0\, Y => \U1/N_266\);
    
    \U1/data_all[233]\ : DFN1E0C0
      port map(D => \U1/N_223\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[233]\);
    
    \U5/data_send_RNO_0[5]\ : MX2C
      port map(A => \U5/N_520\, B => \U5/N_528\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i69_mux\);
    
    \U1/data_all[15]\ : DFN1E0C0
      port map(D => \U1/data_all_3[15]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[15]\);
    
    \U2/parity_check_RNO_15\ : NOR3B
      port map(A => \U2/N_178\, B => \U2/N_173\, C => \U2/N_59_i\, 
        Y => \U2/N_118\);
    
    \U1/data_all_RNO_0[51]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[51]\, Y => 
        \U1/N_2151\);
    
    \U1/data_all_RNO_0[216]\ : AO1C
      port map(A => \data_all[216]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m64_1_i_0_0\);
    
    \U1/data_all_RNO[27]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2255\, C
         => \U1/N_2256\, Y => \U1/N_1792\);
    
    \U1/data_all[56]\ : DFN1E0C0
      port map(D => \U1/N_690\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[56]\);
    
    \U1/data_all[193]\ : DFN1E0C0
      port map(D => \U1/N_96\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[193]\);
    
    \U5/data_send_RNO_10[7]\ : MX2
      port map(A => \U5/N_410\, B => \U5/N_418\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_498\);
    
    \U1/data_all_RNO_0[22]\ : AO1C
      port map(A => \data_all[22]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m147_0_0_i_0\);
    
    \addr_pad[2]/U0/U0\ : IOPAD_TRI
      port map(D => \addr_pad[2]/U0/NET1\, E => 
        \addr_pad[2]/U0/NET2\, PAD => addr(2));
    
    \U5/data_send_RNO_8[6]\ : MX2
      port map(A => \U5/N_377\, B => \U5/N_385\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_481\);
    
    \U2/cnt_RNI05BL9[1]\ : OR3
      port map(A => \U2/N_111\, B => \U2/N_114\, C => 
        \U2/un1_tx_uart27_1_0\, Y => \U2/un1_tx_uart27_4_2\);
    
    \U5/data_send_RNO[7]\ : MX2A
      port map(A => \U5/i58_mux\, B => \U5/N_27_0\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[7]\);
    
    \U5/data_send[0]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[0]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[0]\);
    
    \U1/cnt_daly_RNICDTJ4[8]\ : NOR2B
      port map(A => \U1/m20_m6_0_a2_7\, B => \U1/m20_m6_0_a2_6\, 
        Y => \U1/m20_N_13_mux\);
    
    \U1/data_all[127]\ : DFN1E0C0
      port map(D => \U1/N_70\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[127]\);
    
    \U5/data_send_RNO_1[5]\ : MX2A
      port map(A => \U5/N_116\, B => \U5/N_40_0\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_41_0\);
    
    \U5/data_send_RNO_1[6]\ : MX2A
      port map(A => \U5/N_531\, B => \U5/N_33_0\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_34_0\);
    
    \U2/parity_check_RNO_10\ : XA1A
      port map(A => \data_send[1]\, B => \U2/parity_check_net_1\, 
        C => \U2/parity_check_2_sqmuxa\, Y => \U2/N_119\);
    
    \U1/m107_e_2\ : NOR2B
      port map(A => \data_recive[1]\, B => \data_recive[2]\, Y
         => \U1/m107_e_2_net_1\);
    
    \U0/ce\ : DFN1E0C0
      port map(D => \U0/pr_state[2]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U0/N_138\, Q => ce_c);
    
    \U1/data_all_RNO_0[229]\ : AO1C
      port map(A => \data_all[229]\, B => \U1/N_837_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m89_i_0_0\);
    
    \U1/data_all_RNO_1[230]\ : NOR2
      port map(A => \U1/data_filter[6]_net_1\, B => \U1/N_837\, Y
         => \U1/N_916\);
    
    \U5/cnt_RNI3MVE2[4]\ : NOR3B
      port map(A => \U5/m7_1\, B => \U5/cnt[0]_net_1\, C => 
        \U5/cnt[1]_net_1\, Y => \U5/N_138_mux\);
    
    \U4/pr_state_RNI9BOK1[1]\ : MX2A
      port map(A => \U4/pr_state[1]_net_1\, B => \U4/N_6_0\, S
         => \U4/pr_state[0]_net_1\, Y => \U4/N_7_0\);
    
    \U1/data_all[55]\ : DFN1E0C0
      port map(D => \U1/N_692\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[55]\);
    
    \U2/cnt[6]\ : DFN1C0
      port map(D => \U2/cnt_n6_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[6]_net_1\);
    
    \U0/data_ad_RNO[9]\ : NOR2A
      port map(A => \data_in_c[9]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[9]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I80_un1_Y_0\ : NOR3C
      port map(A => \U1/N245\, B => \U1/N249\, C => \U1/N176\, Y
         => \U1/ADD_14x14_fast_I80_un1_Y_0\);
    
    \data_in_pad[0]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(0), Y => \data_in_pad[0]/U0/NET1\);
    
    \U1/data_all_RNO_0[113]\ : AO1C
      port map(A => \data_all[113]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[113]\);
    
    \U1/data_all_RNO[227]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2159\, C
         => \U1/N_2160\, Y => \U1/N_704\);
    
    \U2/cnt_RNI9CET3[10]\ : OA1
      port map(A => \U2/N_197\, B => \U2/N_192\, C => \U2/N_177\, 
        Y => \U2/un1_tx_uart27_4_1\);
    
    \U5/data_send_RNO_14[1]\ : MX2
      port map(A => \data_all[1]\, B => \data_all[9]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_340\);
    
    \U2/cnt_n6_tz\ : AX1C
      port map(A => \U2/cnt[5]_net_1\, B => \U2/cnt_c4_net_1\, C
         => \U2/cnt[6]_net_1\, Y => \U2/cnt_n6_tz_net_1\);
    
    \U1/data_all_RNO_0[194]\ : AO1C
      port map(A => \data_all[194]\, B => \U1/N_839\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m139_0_i_0\);
    
    \U1/data_all_RNO[21]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m150_i_0_0\, Y => \U1/N_1787\);
    
    \U5/data_send_RNO_17[5]\ : MX2
      port map(A => \data_all[53]\, B => \data_all[61]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_368\);
    
    \U5/data_send_RNO_27[4]\ : MX2
      port map(A => \data_all[212]\, B => \data_all[220]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_447\);
    
    \U1/data_all_RNO[2]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_981\, C
         => \U1/N_982\, Y => \U1/N_2043\);
    
    \U1/data_all_RNO[50]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2153\, C
         => \U1/N_2154\, Y => \U1/N_698\);
    
    \U2/send\ : DFN1E1C0
      port map(D => vld_send, CLK => sys_clk_c, CLR => sys_rest_c, 
        E => \U2/un5_vld_send\, Q => \U2/send_net_1\);
    
    \U1/data_all_RNO_0[117]\ : AO1C
      port map(A => \data_all[117]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[117]\);
    
    \U1/m107_e_3\ : NOR3A
      port map(A => \data_recive[3]\, B => \data_recive[4]\, C
         => \data_recive[7]\, Y => \U1/m107_e_3_net_1\);
    
    \U1/data_all_RNO[121]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[121]\, Y => \U1/N_382\);
    
    \U1/data_all_RNO[234]\ : OA1B
      port map(A => \U1/N_837_0\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[234]\, Y => \U1/N_304\);
    
    \U1/data_all[223]\ : DFN1E0C0
      port map(D => \U1/N_18\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[223]\);
    
    \data_in_pad[5]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(5), Y => \data_in_pad[5]/U0/NET1\);
    
    \U0/conver_ris3\ : DFN1P0
      port map(D => \U0/conver_ris2_i\, CLK => sys_clk_c, PRE => 
        sys_rest_c, Q => \U0/conver_ris3_i_0\);
    
    \U3/cnt_RNIDET01[9]\ : NOR3A
      port map(A => \U3/m106_0\, B => \U3/cnt[4]_net_1\, C => 
        \U3/cnt[9]_net_1\, Y => \U3/m106_5\);
    
    \U2/cnt_RNIUU7J_0[2]\ : NOR2B
      port map(A => \U2/N_131\, B => \U2/N_125\, Y => \U2/N_171\);
    
    \U1/data_all_RNO[223]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_840_0\, C
         => \data_all[223]\, Y => \U1/N_18\);
    
    \U1/data_all[4]\ : DFN1E0C0
      port map(D => \U1/N_255\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[4]\);
    
    \U1/data_all[172]\ : DFN1E0C0
      port map(D => \U1/N_331\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[172]\);
    
    \U0/data_ad_RNO[3]\ : NOR2A
      port map(A => \data_in_c[3]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[3]\);
    
    \U5/data_send_RNO_19[0]\ : MX2
      port map(A => \data_all[80]\, B => \data_all[88]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_379\);
    
    \U4/nx_state_RNO_1[0]\ : NOR2A
      port map(A => \U4/N_23\, B => \U4/pr_state[1]_net_1\, Y => 
        \U4/N_27\);
    
    \U3/receive_over\ : DFN1E0C0
      port map(D => \U3/data_recive31\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U3/receive_over_0_sqmuxa\, Q => 
        receive_over);
    
    \U1/data_all_RNO_1[17]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_836\, Y
         => \U1/N_2276\);
    
    \U1/receive_on_RNIMER81\ : NOR3
      port map(A => receive_on, B => \U1/pr_state[4]_net_1\, C
         => \U1/pr_state[3]_net_1\, Y => \U1/m85_i_0_a3_1\);
    
    \U1/data_all_RNO_0[33]\ : NOR2A
      port map(A => \U1/N_832\, B => \data_all[33]\, Y => 
        \U1/N_2217\);
    
    \U1/cnt_daly[11]\ : DFN1E0C0
      port map(D => \U1/cnt_daly_n11\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => 
        \U1/cnt_daly[11]_net_1\);
    
    \U5/data_send_RNO_10[5]\ : MX2
      port map(A => \U5/N_408\, B => \U5/N_416\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_496\);
    
    \U0/data_ad[8]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[8]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[8]\);
    
    \U5/data_send_RNO_25[7]\ : MX2
      port map(A => \data_all[183]\, B => \data_all[191]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_434\);
    
    \U1/m302_0_i_o2_0_0\ : OR2
      port map(A => \U1/m302_0_i_o2_0_net_1\, B => \U1/N_817\, Y
         => \U1/N_835_0\);
    
    \U1/data_all[89]\ : DFN1E0C0
      port map(D => \U1/N_360\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[89]\);
    
    \U1/data_filter_RNO_0[4]\ : AO1D
      port map(A => \U1/data_filter[6]_net_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, 
        Y => \U1/data_filter_4_i_0_0_0[4]\);
    
    \U1/data_filter[0]\ : DFN1E0C0
      port map(D => \U1/N_61_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[0]_net_1\);
    
    \U1/data_all_RNO[182]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[182]\, Y => \U1/N_405\);
    
    \data_in_pad[4]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(4), Y => \data_in_pad[4]/U0/NET1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I28_Y\ : AO1
      port map(A => \U1/N185\, B => \U1/N189\, C => \U1/N188\, Y
         => \U1/N244\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I25_Y\ : OA1
      port map(A => \U1/data_filter[5]_net_1\, B => \data_ad[5]\, 
        C => \U1/N195\, Y => \U1/N241\);
    
    \U1/data_all_RNO_1[215]\ : NOR2
      port map(A => \U1/data_filter[7]_net_1\, B => \U1/N_840\, Y
         => \U1/N_1022\);
    
    \U1/data_all_RNO_0[104]\ : AO1C
      port map(A => \data_all[104]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[104]\);
    
    \U1/data_all[180]\ : DFN1E0C0
      port map(D => \U1/N_401\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[180]\);
    
    \U5/data_send_RNO_22[0]\ : MX2
      port map(A => \data_all[128]\, B => \data_all[136]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_403\);
    
    \U0/sts_ris\ : DFN1P0
      port map(D => \U0/sts_ris_2\, CLK => sys_clk_c, PRE => 
        sys_rest_c, Q => \U0/sts_ris_i_0\);
    
    \U1/cnt_daly_RNIS0E32[3]\ : OR3B
      port map(A => \U1/cnt_daly[3]_net_1\, B => 
        \U1/cnt_daly[4]_net_1\, C => \U1/N_846\, Y => \U1/N_848\);
    
    \U2/cnt_RNIGILQ4[0]\ : AO1
      port map(A => \U2/tx_uart34_1\, B => \U2/N_194\, C => 
        \U2/tx_uart27\, Y => \U2/un1_tx_uart27_0\);
    
    \U2/cnt_RNI7DUF2_0[10]\ : NOR3C
      port map(A => \U2/N_169\, B => \U2/N_127\, C => \U2/N_181\, 
        Y => \U2/parity_check_1_sqmuxa\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I79_Y_0\ : AO1
      port map(A => \U1/N238\, B => \U1/N235\, C => \U1/N234\, Y
         => \U1/ADD_14x14_fast_I79_Y_0\);
    
    \U5/data_send_RNO_27[6]\ : MX2
      port map(A => \data_all[214]\, B => \data_all[222]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_449\);
    
    \U1/data_all_RNO_0[93]\ : AO1C
      port map(A => \data_all[93]\, B => \U1/N_834_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[93]\);
    
    \U1/data_all_RNO_0[131]\ : AO1C
      port map(A => \data_all[131]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[131]\);
    
    \U4/conver_ris\ : DFN1C0
      port map(D => \U4/conver_ris_2\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U4/conver_ris_net_1\);
    
    \U2/cnt[10]\ : DFN1C0
      port map(D => \U2/cnt_n10_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[10]_net_1\);
    
    \U1/data_all_RNO[96]\ : OA1B
      port map(A => \U1/N_829\, B => \U1/data_filter[0]_net_1\, C
         => \U1/data_all_3_i_0_0_0[96]\, Y => \U1/N_1615\);
    
    \U1/data_all_RNO_0[120]\ : AO1C
      port map(A => \data_all[120]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[120]\);
    
    \U1/data_all[236]\ : DFN1E0C0
      port map(D => \U1/N_30\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[236]\);
    
    \cs_pad/U0/U0\ : IOPAD_TRI
      port map(D => \cs_pad/U0/NET1\, E => \cs_pad/U0/NET2\, PAD
         => cs);
    
    \U1/data_all_RNO_1[209]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_840\, Y
         => \U1/N_1032\);
    
    \U5/data_send_RNO_27[7]\ : MX2
      port map(A => \data_all[215]\, B => \data_all[223]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_450\);
    
    \U1/data_all_RNO_1[217]\ : NOR2
      port map(A => \U1/data_filter[9]_net_1\, B => \U1/N_840\, Y
         => \U1/N_1020\);
    
    \U1/data_all_RNO_0[221]\ : AO1C
      port map(A => \data_all[221]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m57_0_i_0_0\);
    
    \U5/pr_state_RNO[1]\ : NOR3B
      port map(A => send_over, B => \U5/pr_state[0]_net_1\, C => 
        \U5/pr_state[1]_net_1\, Y => \U5/pr_state_RNO[1]_net_1\);
    
    \U2/cnt_RNI8OJ9_0[3]\ : NOR2
      port map(A => \U2/cnt[1]_net_1\, B => \U2/cnt[3]_net_1\, Y
         => \U2/un1_cnt_1\);
    
    \U3/cnt_RNO[0]\ : NOR2A
      port map(A => \U3/recive_net_1\, B => \U3/cnt[0]_net_1\, Y
         => \U3/cnt_4[0]\);
    
    \U2/send_over_RNO\ : OA1
      port map(A => \U2/tx_uart38\, B => \U2/un1_cnt\, C => 
        \U2/send_net_1\, Y => \U2/N_198\);
    
    \U1/data_all_RNO[205]\ : OA1B
      port map(A => \U1/N_839\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m106_i_0_0\, Y => \U1/N_213\);
    
    \U1/data_filter_RNO[0]\ : NOR3
      port map(A => \U1/N_906\, B => \U1/pr_state_0[7]_net_1\, C
         => \U1/N_905\, Y => \U1/N_61_0\);
    
    \U1/data_all_RNO[19]\ : OA1B
      port map(A => \U1/N_836_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/m156_0_i_0_0\, Y => \U1/N_1785\);
    
    \U2/cnt_RNIMDDJ[11]\ : NOR2A
      port map(A => \U2/cnt[11]_net_1\, B => \U2/cnt[0]_net_1\, Y
         => \U2/tx_uart37_0\);
    
    \U3/un7_cnt_1_I_5\ : XOR2
      port map(A => \U3/cnt[0]_net_1\, B => \U3/cnt[1]_net_1\, Y
         => \U3/I_5\);
    
    \U1/data_all_RNO_0[17]\ : NOR2A
      port map(A => \U1/N_836\, B => \data_all[17]\, Y => 
        \U1/N_2275\);
    
    \U2/cnt_RNI7DUF2[0]\ : NOR2B
      port map(A => \U2/N_194\, B => \U2/N_174\, Y => 
        \U2/parity_check_7_sqmuxa\);
    
    \U1/data_all_RNO[108]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[108]\, Y => \U1/N_1611\);
    
    \U1/conver_RNO\ : NOR3
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/pr_state[6]_net_1\, C => \U1/pr_state[7]_net_1\, Y
         => \U1/N_1095\);
    
    \U5/data_send_RNO_12[5]\ : MX2
      port map(A => \U5/N_440\, B => \U5/N_448\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_512\);
    
    \U1/data_all[231]\ : DFN1E0C0
      port map(D => \U1/N_32\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[231]\);
    
    \U1/data_all[133]\ : DFN1E0C0
      port map(D => \U1/N_1836\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[133]\);
    
    \U5/data_send_RNO_7[5]\ : MX2
      port map(A => \U5/N_360\, B => \U5/N_368\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_472\);
    
    \U5/data_send_RNO_23[1]\ : MX2
      port map(A => \data_all[145]\, B => \data_all[153]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_412\);
    
    \U1/data_all[190]\ : DFN1E0C0
      port map(D => \U1/N_53\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[190]\);
    
    \U0/pr_state_RNO_0[0]\ : OA1C
      port map(A => \U0/pr_state[5]_net_1\, B => 
        \U0/conver_ris_i_0\, C => \U0/pr_state[0]_net_1\, Y => 
        \U0/N_143\);
    
    \U5/data_send_RNO_2[2]\ : MX2
      port map(A => \U5/N_461\, B => \U5/N_469\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_517\);
    
    \U1/data_all_RNO_0[34]\ : AO1C
      port map(A => \data_all[34]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m292_i_0_0\);
    
    \U1/data_all_RNO_0[43]\ : NOR2A
      port map(A => \U1/N_832\, B => \data_all[43]\, Y => 
        \U1/N_2197\);
    
    \U1/data_all_RNO_0[185]\ : AO1C
      port map(A => \data_all[185]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[185]\);
    
    \U1/data_all_RNO[236]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_983\, C
         => \U1/N_984\, Y => \U1/N_30\);
    
    \U1/data_all_RNO_1[57]\ : NOR2
      port map(A => \U1/data_filter[9]_net_1\, B => \U1/N_831\, Y
         => \U1/N_2144\);
    
    \U0/cnt_rc_n0\ : NOR2
      port map(A => \U0/cnt_rc[0]_net_1\, B => 
        \U0/pr_state[4]_net_1\, Y => \U0/N_164\);
    
    \U1/data_all[19]\ : DFN1E0C0
      port map(D => \U1/N_1785\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[19]\);
    
    \U1/data_all[155]\ : DFN1E0C0
      port map(D => \U1/N_1801\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[155]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I99_Y\ : AX1D
      port map(A => \U1/I62_un1_Y\, B => 
        \U1/ADD_14x14_fast_I78_Y_1\, C => 
        \U1/ADD_14x14_fast_I99_Y_0\, Y => 
        \U1/un2_data_filter[11]\);
    
    \U1/un14_data_all_I_11\ : NOR2
      port map(A => \U1/DWACT_FDEC_E[0]\, B => \addr_c[3]\, Y => 
        \U1/OVER\);
    
    \U5/data_send_RNO_7[2]\ : MX2
      port map(A => \U5/N_357\, B => \U5/N_365\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_469\);
    
    \U3/cnt_RNI1TAQ1[4]\ : NOR3C
      port map(A => \U3/m11_3\, B => \U3/m11_2\, C => \U3/m11_6\, 
        Y => \U3/m11_9\);
    
    \U0/pr_state_RNO[3]\ : AO1
      port map(A => \U0/sts_ris_i_0\, B => \U0/pr_state[3]_net_1\, 
        C => \U0/pr_state[4]_net_1\, Y => \U0/pr_state_ns[2]\);
    
    \U5/data_send_RNO_13[0]\ : NOR2A
      port map(A => \U5/N_451\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_74\);
    
    \U1/data_all_RNO_1[49]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_831\, Y
         => \U1/N_2156\);
    
    \U2/cnt_RNIH1K9_0[8]\ : NOR2A
      port map(A => \U2/cnt[8]_net_1\, B => \U2/cnt[5]_net_1\, Y
         => \U2/un1_cnt_3\);
    
    \U1/cnt_daly_RNO_1[8]\ : OA1C
      port map(A => \U1/cnt_daly[7]_net_1\, B => \U1/N_850\, C
         => \U1/cnt_daly[8]_net_1\, Y => \U1/N_2303\);
    
    \U5/data_send_RNO_2[3]\ : MX2
      port map(A => \U5/N_462\, B => \U5/N_470\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_518\);
    
    \U2/cnt_RNI8PAD2[1]\ : NOR3C
      port map(A => \U2/tx_uart27_0_a2_2\, B => 
        \U2/tx_uart27_0_a2_1\, C => \U2/tx_uart27_0_a2_3\, Y => 
        \U2/tx_uart27\);
    
    \U1/data_all[226]\ : DFN1E0C0
      port map(D => \U1/N_706\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[226]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I48_Y\ : AO1
      port map(A => \U1/N244\, B => \U1/N241\, C => \U1/N240\, Y
         => \U1/N267\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I45_Y\ : NOR2B
      port map(A => \U1/N241\, B => \U1/N237\, Y => \U1/N264\);
    
    \U0/cnt_rc_n2\ : XA1C
      port map(A => \U0/N_130\, B => \U0/cnt_rc[2]_net_1\, C => 
        \U0/pr_state[4]_net_1\, Y => \U0/cnt_rc_n2_net_1\);
    
    \U5/data_send_RNO_7[3]\ : MX2
      port map(A => \U5/N_358\, B => \U5/N_366\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_470\);
    
    \U5/data_send_RNO_21[6]\ : MX2
      port map(A => \data_all[118]\, B => \data_all[126]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_401\);
    
    \U3/data_recive_RNO_2[0]\ : NOR3A
      port map(A => \U3/m36_1\, B => \U3/cnt[10]_net_1\, C => 
        \U3/cnt[7]_net_1\, Y => \U3/m62_5\);
    
    \U1/data_all[59]\ : DFN1E0C0
      port map(D => \U1/N_680\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[59]\);
    
    \U3/data_recive_RNO_1[0]\ : NOR3C
      port map(A => \U3/m62_5\, B => \U3/N_39\, C => \U3/m62_6\, 
        Y => \U3/data_recive23\);
    
    \U1/data_all_RNO_0[66]\ : AO1C
      port map(A => \data_all[66]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m246_i_0_0\);
    
    \U1/data_all_RNO_0[50]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[50]\, Y => 
        \U1/N_2153\);
    
    \U5/data_send_RNO_26[0]\ : MX2
      port map(A => \data_all[192]\, B => \data_all[200]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_435\);
    
    \U1/data_all[64]\ : DFN1E0C0
      port map(D => \U1/N_163\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[64]\);
    
    \U1/cnt_daly[7]\ : DFN1E0C0
      port map(D => \U1/N_808\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[7]_net_1\);
    
    \U5/data_send_RNO_15[6]\ : MX2
      port map(A => \data_all[22]\, B => \data_all[30]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_353\);
    
    \U3/data_recive_RNO[6]\ : MX2
      port map(A => \U3/m81_0\, B => rx_uart_c, S => 
        \U3/data_recive29\, Y => \U3/data_recive_12[6]\);
    
    \U1/data_all_RNO_0[69]\ : AO1C
      port map(A => \data_all[69]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m237_i_0_0\);
    
    \U1/cnt_daly_RNO[2]\ : XA1C
      port map(A => \U1/cnt_daly[2]_net_1\, B => \U1/N_845\, C
         => \U1/pr_state[7]_net_1\, Y => \U1/N_798\);
    
    \U5/data_send_RNO_5[4]\ : MX2
      port map(A => \U5/N_511\, B => \U5/N_46_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_47_0\);
    
    \U5/data_send_RNO_10[0]\ : MX2
      port map(A => \U5/N_403\, B => \U5/N_411\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_491\);
    
    \U1/pr_state_RNO[0]\ : NOR3
      port map(A => \U1/N_864\, B => \U1/N_866\, C => \U1/N_865\, 
        Y => \U1/pr_state_RNO[0]_net_1\);
    
    \U1/data_all_RNO_1[20]\ : NOR2
      port map(A => \U1/data_filter[4]_net_1\, B => \U1/N_836\, Y
         => \U1/N_2270\);
    
    \U1/data_filter_RNO_0[2]\ : AO1D
      port map(A => \U1/data_filter[4]_net_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, 
        Y => \U1/data_filter_4_i_0_0_0[2]\);
    
    \U1/data_all[221]\ : DFN1E0C0
      port map(D => \U1/N_1780\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[221]\);
    
    \U1/data_all[123]\ : DFN1E0C0
      port map(D => \U1/N_386\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[123]\);
    
    \U1/data_all_RNO_1[3]\ : NOR2
      port map(A => \U1/data_filter[3]_net_1\, B => \U1/N_835\, Y
         => \U1/N_1097\);
    
    \U2/cnt_RNIEM1T[5]\ : NOR3A
      port map(A => \U2/tx_uart37_6\, B => \U2/cnt[7]_net_1\, C
         => \U2/cnt[5]_net_1\, Y => \U2/tx_uart38_1\);
    
    \U1/m253_i_0_o2_0_0\ : OR2
      port map(A => \U1/m253_i_0_o2_0_net_1\, B => \U1/N_817\, Y
         => \U1/N_832_0\);
    
    \U1/data_all[60]\ : DFN1E0C0
      port map(D => \U1/N_31\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[60]\);
    
    \U1/data_all_RNO[37]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m283_i_0_0\, Y => \U1/N_1810\);
    
    \U1/data_all_RNO[169]\ : OA1B
      port map(A => \U1/N_838\, B => \U1/data_filter[9]_net_1\, C
         => \U1/m167_i_0_0\, Y => \U1/N_325\);
    
    \U5/data_send_RNO_15[3]\ : MX2
      port map(A => \data_all[19]\, B => \data_all[27]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_350\);
    
    \U1/data_all_RNO_1[55]\ : NOR2
      port map(A => \U1/data_filter[7]_net_1\, B => \U1/N_831\, Y
         => \U1/N_2148\);
    
    \U1/data_all_RNO_0[189]\ : AO1C
      port map(A => \data_all[189]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[189]\);
    
    \U1/data_all_RNO_0[26]\ : AO1C
      port map(A => \data_all[26]\, B => \U1/N_836\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m135_0_i_0_0\);
    
    \U1/data_all[218]\ : DFN1E0C0
      port map(D => \U1/N_1778\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[218]\);
    
    \U1/data_all_RNO_0[186]\ : NOR2A
      port map(A => \U1/N_844\, B => \data_all[186]\, Y => 
        \U1/N_2081\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I68_un1_Y\ : NOR3C
      port map(A => \U1/N243\, B => \U1/N239\, C => \U1/N273\, Y
         => \U1/I68_un1_Y\);
    
    \U1/data_all_RNO_0[29]\ : AO1C
      port map(A => \data_all[29]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m125_0_0_i_0\);
    
    \U1/data_all_RNO_0[182]\ : AO1C
      port map(A => \data_all[182]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[182]\);
    
    \U2/cnt_RNICSJ9_1[2]\ : NOR2
      port map(A => \U2/cnt[2]_net_1\, B => \U2/cnt[6]_net_1\, Y
         => \U2/tx_uart36_5\);
    
    \U1/data_all_RNO_0[44]\ : AO1C
      port map(A => \data_all[44]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m261_i_0_0\);
    
    \U1/cnt_daly_RNIL3VQ[1]\ : OR2B
      port map(A => \U1/cnt_daly[1]_net_1\, B => 
        \U1/cnt_daly[0]_net_1\, Y => \U1/N_845\);
    
    \U1/receive_flag_RNO\ : AO1
      port map(A => \U1/m112_i_0_a3_0\, B => \U1/N_139\, C => 
        addr_over, Y => \U1/N_263\);
    
    \U1/data_all_3_i_o3_0_o2_0_o2_0[143]\ : OR3B
      port map(A => \addr_c_0[0]\, B => \U1/I_9_0\, C => 
        \U1/I_5_0\, Y => \U1/m103_i_o2_0_o2_0_net_1\);
    
    \U1/cnt_daly_RNI1NE81[1]\ : OR3C
      port map(A => \U1/cnt_daly[0]_net_1\, B => 
        \U1/cnt_daly[1]_net_1\, C => \U1/cnt_daly[2]_net_1\, Y
         => \U1/N_846\);
    
    \U1/data_all_RNO[132]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[132]\, Y => \U1/N_245\);
    
    \U1/data_all[66]\ : DFN1E0C0
      port map(D => \U1/N_167\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[66]\);
    
    \U3/data_recive_RNO_2[1]\ : NOR3A
      port map(A => \U3/cnt[3]_net_1\, B => \U3/cnt[5]_net_1\, C
         => \U3/cnt[10]_net_1\, Y => \U3/m27_2\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I76_Y\ : AO1
      port map(A => \U1/ADD_14x14_fast_I76_un1_Y_0\, B => 
        \U1/N332\, C => \U1/ADD_14x14_fast_I76_Y_1\, Y => 
        \U1/N313\);
    
    \U1/data_all_RNO_0[188]\ : AO1C
      port map(A => \data_all[188]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[188]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I77_Y_2\ : AO1
      port map(A => \U1/N258\, B => \U1/N265\, C => 
        \U1/ADD_14x14_fast_I77_Y_1\, Y => 
        \U1/ADD_14x14_fast_I77_Y_2\);
    
    \U1/data_all_RNO[20]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2269\, C
         => \U1/N_2270\, Y => \U1/N_1786\);
    
    \U1/data_all_3_0_0_i_o2[220]\ : OR2
      port map(A => \U1/m79_0_i_i_o2_0_net_1\, B => \U1/N_818\, Y
         => \U1/N_840\);
    
    \U1/data_all[171]\ : DFN1E0C0
      port map(D => \U1/N_329\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[171]\);
    
    \U0/cnt_rc[2]\ : DFN1E0C0
      port map(D => \U0/cnt_rc_n2_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U0/N_135\, Q => 
        \U0/cnt_rc[2]_net_1\);
    
    \U3/data_recive_RNO_3[2]\ : NOR3C
      port map(A => \U3/cnt[7]_net_1\, B => \U3/cnt[2]_net_1\, C
         => \U3/m11_3\, Y => \U3/m70_4\);
    
    \U1/data_all_RNO[185]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[185]\, Y => \U1/N_411\);
    
    \U1/data_all[93]\ : DFN1E0C0
      port map(D => \U1/N_1776\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[93]\);
    
    \U5/data_send_RNO_14[2]\ : MX2
      port map(A => \data_all[2]\, B => \data_all[10]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_341\);
    
    \U5/data_send_RNO_11[1]\ : MX2
      port map(A => \U5/N_420\, B => \U5/N_428\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_500\);
    
    \U2/tx_uart_RNO_0\ : OA1A
      port map(A => \U2/un1_tx_uart27\, B => \U2/tx_uart38\, C
         => \U2/send_net_1\, Y => \U2/tx_uart_11_sqmuxa\);
    
    \U1/data_all_RNO[6]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[6]\, Y => \U1/N_250\);
    
    \data_in_pad[10]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(10), Y => \data_in_pad[10]/U0/NET1\);
    
    \U1/data_all_RNO[31]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_836\, C
         => \data_all[31]\, Y => \U1/data_all_3[31]\);
    
    \U5/data_send_RNO_13[7]\ : NOR2A
      port map(A => \U5/N_458\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_25_0\);
    
    \U3/cnt[11]\ : DFN1C0
      port map(D => \U3/cnt_4[11]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U3/cnt[11]_net_1\);
    
    \U2/tx_uart_RNO_5\ : NOR2B
      port map(A => \U2/parity_check_3_sqmuxa\, B => 
        \data_send[2]\, Y => \U2/data_send_m[2]\);
    
    \U1/un14_data_all_I_10\ : OR3
      port map(A => \addr_c[0]\, B => \addr_c[1]\, C => 
        \addr_c[2]\, Y => \U1/DWACT_FDEC_E[0]\);
    
    \U1/data_all_RNO[192]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/m145_i_0_0\, Y => \U1/N_197\);
    
    \U1/data_all[65]\ : DFN1E0C0
      port map(D => \U1/N_165\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[65]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I34_Y\ : AO1
      port map(A => \U1/N180\, B => \U1/N176\, C => \U1/N179\, Y
         => \U1/N250\);
    
    \U1/data_all_RNO[179]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[179]\, Y => \U1/N_399\);
    
    \U1/data_all_RNO[16]\ : OA1B
      port map(A => \U1/N_836\, B => \U1/data_filter[0]_net_1\, C
         => \U1/m163_0_i_0_0\, Y => \U1/N_1782\);
    
    \U5/data_send_RNO_2[6]\ : MX2
      port map(A => \U5/N_465\, B => \U5/N_473\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_521\);
    
    \U2/tx_uart_RNO_11\ : NOR2B
      port map(A => \U2/parity_check_7_sqmuxa\, B => 
        \data_send[6]\, Y => \U2/data_send_m[6]\);
    
    \U5/data_send_RNO_20[3]\ : MX2
      port map(A => \data_all[99]\, B => \data_all[107]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_390\);
    
    \U1/data_all_RNO[207]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[207]\, 
        C => \U1/N_839\, Y => \U1/N_158\);
    
    \U1/data_all[146]\ : DFN1E0C0
      port map(D => \U1/N_1796\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[146]\);
    
    \U1/data_all_RNO[159]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_842_0\, C
         => \data_all[159]\, Y => \U1/data_all_3[159]\);
    
    \data_in_pad[7]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(7), Y => \data_in_pad[7]/U0/NET1\);
    
    \U1/data_all[166]\ : DFN1E0C0
      port map(D => \U1/N_319\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[166]\);
    
    \U3/data_recive_RNO[0]\ : MX2
      port map(A => \U3/m93_0\, B => rx_uart_c, S => 
        \U3/data_recive23\, Y => \U3/data_recive_12[0]\);
    
    \U2/cnt_RNIH1K9_1[8]\ : NOR2A
      port map(A => \U2/cnt[5]_net_1\, B => \U2/cnt[8]_net_1\, Y
         => \U2/un1_tx_uart27_3_0_a2_3_0\);
    
    \U1/data_all[208]\ : DFN1E0C0
      port map(D => \U1/N_196\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[208]\);
    
    \U1/data_all_RNO[101]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[101]\, Y => \U1/N_56\);
    
    \U1/pr_state_RNIU1MS[0]\ : OR2
      port map(A => \U1/pr_state[0]_net_1\, B => 
        \U1/pr_state[2]_net_1\, Y => \U1/N_854\);
    
    \U1/data_all_3_i_0_0_o2_0[190]\ : OR2
      port map(A => \U1/data_all_3_i_0_0_o2_1[190]_net_1\, B => 
        \U1/N_817\, Y => \U1/N_844_0\);
    
    \U2/tx_uart_RNO_10\ : AO1B
      port map(A => \U2/tx_uart37_8\, B => \U2/tx_uart37_7\, C
         => \U2/send_net_1\, Y => \U2/tx_uart_11_iv_0\);
    
    \U1/data_all[130]\ : DFN1E0C0
      port map(D => \U1/N_107\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[130]\);
    
    \U3/cnt_RNIFGT01[6]\ : NOR3C
      port map(A => \U3/cnt[7]_net_1\, B => \U3/cnt[6]_net_1\, C
         => \U3/m11_3\, Y => \U3/m106_6\);
    
    \data_in_pad[11]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(11), Y => \data_in_pad[11]/U0/NET1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I5_G0N\ : NOR2B
      port map(A => \data_ad[5]\, B => \U1/data_filter[5]_net_1\, 
        Y => \U1/N191\);
    
    \U3/cnt_RNIKFN33[1]\ : NOR2B
      port map(A => \U3/m11_9\, B => \U3/m11_8\, Y => 
        \U3/data_recive31\);
    
    \U5/data_send_RNO_13[4]\ : NOR2A
      port map(A => \U5/N_455\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_46_0\);
    
    \U2/cnt_RNI8OJ9[3]\ : NOR2B
      port map(A => \U2/cnt[3]_net_1\, B => \U2/cnt[1]_net_1\, Y
         => \U2/tx_uart37_1\);
    
    \U1/data_all_RNO[203]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[11]_net_1\, 
        C => \U1/m112_0_0_i_0\, Y => \U1/N_75\);
    
    \U3/data_recive_RNO_2[4]\ : NOR3B
      port map(A => \U3/cnt[0]_net_1\, B => \U3/m22_0\, C => 
        \U3/cnt[8]_net_1\, Y => \U3/m53_3\);
    
    \U2/cnt_RNIDTJ9[3]\ : NOR2A
      port map(A => \U2/cnt[6]_net_1\, B => \U2/cnt[3]_net_1\, Y
         => \U2/tx_uart38_10_1\);
    
    \U2/tx_uart_RNO_9\ : NOR3C
      port map(A => \U2/N_178\, B => \U2/N_173\, C => 
        \data_send[3]\, Y => \U2/data_send_m[3]\);
    
    \U5/data_send_RNO_13[3]\ : NOR2A
      port map(A => \U5/N_454\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_53_0\);
    
    \U1/data_all[115]\ : DFN1E0C0
      port map(D => \U1/N_370\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[115]\);
    
    \U1/data_all_RNO_0[101]\ : AO1C
      port map(A => \data_all[101]\, B => \U1/N_829\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[101]\);
    
    \U0/data_ad[1]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[1]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[1]\);
    
    \U1/data_all_RNO_0[215]\ : NOR2A
      port map(A => \U1/N_840\, B => \data_all[215]\, Y => 
        \U1/N_1021\);
    
    \U5/data_send_RNO_8[5]\ : MX2
      port map(A => \U5/N_376\, B => \U5/N_384\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_480\);
    
    \U5/data_send_RNO_20[1]\ : MX2
      port map(A => \data_all[97]\, B => \data_all[105]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_388\);
    
    \U2/parity_check_RNO_6\ : XA1A
      port map(A => \data_send[5]\, B => \U2/parity_check_net_1\, 
        C => \U2/parity_check_6_sqmuxa\, Y => \U2/N_120\);
    
    \sys_clk_pad/U0/U1\ : CLKIO
      port map(A => \sys_clk_pad/U0/NET1\, Y => sys_clk_c);
    
    \U2/tx_uart_RNO_3\ : OR3
      port map(A => \U2/data_send_m[7]\, B => 
        \U2/tx_uart_11_iv_1\, C => \U2/tx_uart_11_iv_3\, Y => 
        \U2/tx_uart_11_iv_7\);
    
    \U1/cnt_daly_RNIBNTG2[2]\ : NOR3B
      port map(A => \U1/m20_m6_0_a2_2\, B => \U1/m20_m6_0_a2_1\, 
        C => \U1/N_845\, Y => \U1/m20_m6_0_a2_7\);
    
    \U5/data_send_RNO_13[5]\ : NOR2A
      port map(A => \U5/N_456\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_39_0\);
    
    \U2/cnt[7]\ : DFN1C0
      port map(D => \U2/cnt_n7_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[7]_net_1\);
    
    \U1/data_all_RNO_0[88]\ : AO1C
      port map(A => \data_all[88]\, B => \U1/N_834_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[88]\);
    
    \U1/data_all[98]\ : DFN1E0C0
      port map(D => \U1/N_1613\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[98]\);
    
    \U1/data_all[44]\ : DFN1E0C0
      port map(D => \U1/N_290\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[44]\);
    
    \U1/data_all[152]\ : DFN1E0C0
      port map(D => \U1/N_1798\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[152]\);
    
    \U3/cnt_RNID9UG[7]\ : NOR2
      port map(A => \U3/cnt[7]_net_1\, B => \U3/cnt[0]_net_1\, Y
         => \U3/m17_1\);
    
    \U2/cnt_RNI5MRS_0[0]\ : NOR3C
      port map(A => \U2/N_166\, B => \U2/N_124\, C => \U2/N_126\, 
        Y => \U2/N_169\);
    
    \U1/data_all_RNO[44]\ : OA1B
      port map(A => \U1/N_832_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/m261_i_0_0\, Y => \U1/N_290\);
    
    \U1/data_all_RNO[187]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2079\, C
         => \U1/N_2080\, Y => \U1/N_415\);
    
    \addr_pad[3]/U0/U1\ : IOTRI_OB_EB
      port map(D => \addr_c[3]\, E => \VCC\, DOUT => 
        \addr_pad[3]/U0/NET1\, EOUT => \addr_pad[3]/U0/NET2\);
    
    \U5/data_send_RNO_21[4]\ : MX2
      port map(A => \data_all[116]\, B => \data_all[124]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_399\);
    
    \U1/data_all_RNO[126]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[126]\, 
        C => \U1/N_830\, Y => \U1/N_72\);
    
    \U3/rx_down\ : DFN1C0
      port map(D => \U3/rx_down_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/rx_down_net_1\);
    
    \U1/cnt_n1\ : XA1B
      port map(A => \U1/cnt[1]_net_1\, B => \U1/cnt[0]_net_1\, C
         => \U1/pr_state_0[7]_net_1\, Y => \U1/cnt_n1_net_1\);
    
    \U1/data_all[40]\ : DFN1E0C0
      port map(D => \U1/N_266\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[40]\);
    
    \U1/data_all[120]\ : DFN1E0C0
      port map(D => \U1/N_380\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[120]\);
    
    \U1/data_all_RNO_0[3]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[3]\, Y => 
        \U1/N_1096\);
    
    \U1/data_all[149]\ : DFN1E0C0
      port map(D => \U1/N_1797\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[149]\);
    
    \U3/cnt_RNI0URH1[7]\ : NOR3C
      port map(A => \U3/m41_0\, B => \U3/cnt[7]_net_1\, C => 
        \U3/N_39\, Y => \U3/N_120_mux\);
    
    \U1/data_all_RNO_0[53]\ : AO1C
      port map(A => \data_all[53]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[53]\);
    
    \U1/data_all_RNO_0[81]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[81]\, Y => 
        \U1/N_2073\);
    
    \U1/data_all_RNO_0[124]\ : AO1C
      port map(A => \data_all[124]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[124]\);
    
    \U1/data_all_3_0_0_i_o2_0[220]\ : OR2
      port map(A => \U1/m79_0_i_i_o2_0_net_1\, B => \U1/N_818\, Y
         => \U1/N_840_0\);
    
    \U5/data_send_RNO_3[6]\ : MX2
      port map(A => \U5/N_481\, B => \U5/N_489\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_529\);
    
    \U1/pr_state_0[7]\ : DFN1P0
      port map(D => \U1/pr_state_RNICDI39[1]_net_1\, CLK => 
        sys_clk_c, PRE => sys_rest_c, Q => 
        \U1/pr_state_0[7]_net_1\);
    
    \U1/data_all[169]\ : DFN1E0C0
      port map(D => \U1/N_325\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[169]\);
    
    \U5/data_send_RNO_8[7]\ : MX2
      port map(A => \U5/N_378\, B => \U5/N_386\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_482\);
    
    \U1/cnt_daly[6]\ : DFN1E0C0
      port map(D => \U1/N_806\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[6]_net_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I19_Y\ : NOR2B
      port map(A => \U1/N204\, B => \U1/N201\, Y => \U1/N235\);
    
    \U1/data_all[46]\ : DFN1E0C0
      port map(D => \U1/data_all_3[46]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[46]\);
    
    \U1/data_all[105]\ : DFN1E0C0
      port map(D => \U1/N_1612\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[105]\);
    
    \U2/parity_check_RNO_14\ : XOR2
      port map(A => \data_send[6]\, B => \U2/parity_check_net_1\, 
        Y => \U2/N_55_i\);
    
    \U5/data_send_RNO_11[7]\ : MX2
      port map(A => \U5/N_426\, B => \U5/N_434\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_506\);
    
    \U0/data_ad[0]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[0]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[0]\);
    
    \U5/data_send_RNO_10[4]\ : MX2
      port map(A => \U5/N_407\, B => \U5/N_415\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_495\);
    
    \U5/data_send_RNO_8[2]\ : MX2
      port map(A => \U5/N_373\, B => \U5/N_381\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_477\);
    
    \U1/data_all_RNO[54]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[54]\, Y => \U1/N_43\);
    
    \U1/data_all_RNO[135]\ : OA1B
      port map(A => \U1/N_841\, B => \U1/data_filter[7]_net_1\, C
         => \U1/m202_0_i_0\, Y => \U1/N_105\);
    
    \U1/data_all[92]\ : DFN1E0C0
      port map(D => \U1/N_199\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[92]\);
    
    \U1/data_all_RNO[222]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_840_0\, C
         => \data_all[222]\, Y => \U1/N_1781\);
    
    \U0/cnt_rc_RNIJ0US[2]\ : AND3B
      port map(A => \U0/cnt_rc[2]_net_1\, B => 
        \U0/cnt_rc[0]_net_1\, C => \U0/pr_state_ns_a4_2[1]\, Y
         => \U0/pr_state_ns[1]\);
    
    \U3/data_recive_RNO[7]\ : MX2
      port map(A => \U3/m72_0\, B => rx_uart_c, S => 
        \U3/data_recive30\, Y => \U3/data_recive_12[7]\);
    
    \U2/cnt[2]\ : DFN1C0
      port map(D => \U2/cnt_n2_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[2]_net_1\);
    
    \U1/data_all[178]\ : DFN1E0C0
      port map(D => \U1/N_397\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[178]\);
    
    \U5/send_whole_over\ : DFN1E1C0
      port map(D => \U5/pr_state[1]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/un1_pr_state_1\, Q => 
        send_whole_over);
    
    \U1/data_all[45]\ : DFN1E0C0
      port map(D => \U1/N_296\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[45]\);
    
    \U5/data_send_RNO_3[5]\ : MX2
      port map(A => \U5/N_480\, B => \U5/N_488\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_528\);
    
    \U1/data_all[235]\ : DFN1E0C0
      port map(D => \U1/N_225\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[235]\);
    
    \U1/data_all_RNO_0[180]\ : AO1C
      port map(A => \data_all[180]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[180]\);
    
    \U3/cnt_RNICFEO[11]\ : NOR3A
      port map(A => \U3/cnt[11]_net_1\, B => \U3/cnt[9]_net_1\, C
         => \U3/cnt[8]_net_1\, Y => \U3/m11_4\);
    
    \U5/data_send_RNO_4[3]\ : MX2C
      port map(A => \U5/N_494\, B => \U5/N_502\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_534\);
    
    \U1/data_all_RNO[123]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[11]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[123]\, Y => \U1/N_386\);
    
    \U1/data_all_RNO[120]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[120]\, Y => \U1/N_380\);
    
    \U0/cnt_rc_c1_i\ : OR2B
      port map(A => \U0/cnt_rc[1]_net_1\, B => 
        \U0/cnt_rc[0]_net_1\, Y => \U0/N_130\);
    
    \U1/data_all_RNO[195]\ : OA1B
      port map(A => \U1/N_839\, B => \U1/data_filter[3]_net_1\, C
         => \U1/m136_i_0_0\, Y => \U1/N_201\);
    
    \U2/cnt_RNI7NJ9[0]\ : NOR2B
      port map(A => \U2/cnt[0]_net_1\, B => \U2/cnt[3]_net_1\, Y
         => \U2/N_126\);
    
    \U3/un7_cnt_1_I_10\ : AND3
      port map(A => \U3/cnt[0]_net_1\, B => \U3/cnt[1]_net_1\, C
         => \U3/cnt[2]_net_1\, Y => \U3/DWACT_FINC_E[0]\);
    
    \U1/cnt_daly_RNO_0[9]\ : NOR3B
      port map(A => \U1/m24_m4_e_4\, B => \U1/m24_m4_e_3\, C => 
        \U1/N_845\, Y => \U1/m24_N_11_mux\);
    
    \U2/cnt_RNIHP1T[8]\ : NOR3A
      port map(A => \U2/tx_uart37_6\, B => \U2/cnt[7]_net_1\, C
         => \U2/cnt[8]_net_1\, Y => \U2/tx_uart37_7\);
    
    \U1/data_all[69]\ : DFN1E0C0
      port map(D => \U1/N_173\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[69]\);
    
    \U5/data_send_RNO_10[2]\ : MX2
      port map(A => \U5/N_405\, B => \U5/N_413\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_493\);
    
    \U1/data_all_RNO_0[54]\ : AO1C
      port map(A => \data_all[54]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[54]\);
    
    \U1/data_all_RNO[78]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_833\, C
         => \data_all[78]\, Y => \U1/data_all_3[78]\);
    
    \U4/addr[0]\ : DFN1E0C0
      port map(D => \U4/N_20\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U4/N_7_0\, Q => \addr_c[0]\);
    
    \U1/pr_state_RNI02BE[2]\ : CLKINT
      port map(A => \U1/pr_state_0[2]\, Y => 
        \U1/pr_state[2]_net_1\);
    
    \U0/conver_ris\ : DFN1P0
      port map(D => \U0/conver_ris_1\, CLK => sys_clk_c, PRE => 
        sys_rest_c, Q => \U0/conver_ris_i_0\);
    
    \U3/un7_cnt_1_I_30\ : AND3
      port map(A => \U3/DWACT_FINC_E[0]\, B => 
        \U3/DWACT_FINC_E[2]\, C => \U3/DWACT_FINC_E[5]\, Y => 
        \U3/DWACT_FINC_E[6]\);
    
    \U1/cnt_daly_RNO_0[4]\ : OA1C
      port map(A => \U1/cnt_daly[3]_net_1\, B => \U1/N_846\, C
         => \U1/cnt_daly[4]_net_1\, Y => \U1/N_2299\);
    
    \U1/data_all[91]\ : DFN1E0C0
      port map(D => \U1/N_362\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[91]\);
    
    \U1/data_all_RNO_0[165]\ : AO1C
      port map(A => \data_all[165]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m179_i_0_0\);
    
    \U3/idle_recive_RNO\ : INV
      port map(A => \U3/recive_net_1\, Y => \U3/recive_i\);
    
    \U1/data_all[97]\ : DFN1E0C0
      port map(D => \U1/N_1614\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[97]\);
    
    \U1/pr_state_RNO_0[0]\ : OA1B
      port map(A => \U1/N_856\, B => \U1/N_860\, C => \U1/N_854\, 
        Y => \U1/N_864\);
    
    \U1/data_all_RNO_0[32]\ : AO1C
      port map(A => \data_all[32]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m298_i_0_0\);
    
    \U1/data_all_RNO[30]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_836\, C
         => \data_all[30]\, Y => \U1/data_all_3[30]\);
    
    \U1/data_all[225]\ : DFN1E0C0
      port map(D => \U1/N_708\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[225]\);
    
    \U0/cnt_rc_8\ : NOR2A
      port map(A => \U0/cnt_rc[3]_net_1\, B => 
        \U0/pr_state[4]_net_1\, Y => \U0/N_59\);
    
    \U5/data_send_RNO_3[7]\ : MX2C
      port map(A => \U5/N_482\, B => \U5/N_490\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_538\);
    
    \U1/data_all_RNO_1[81]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_834\, Y
         => \U1/N_1050\);
    
    \U5/data_send_RNO_28[1]\ : MX2
      port map(A => \data_all[225]\, B => \data_all[233]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_452\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I98_Y\ : XOR3
      port map(A => \U1/data_filter[10]_net_1\, B => 
        \data_ad[10]\, C => \U1/N319\, Y => 
        \U1/un2_data_filter[10]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I95_Y\ : XOR3
      port map(A => \U1/data_filter[7]_net_1\, B => \data_ad[7]\, 
        C => \U1/N326\, Y => \U1/un2_data_filter[7]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I39_Y\ : NOR2B
      port map(A => \U1/N231\, B => \U1/N235\, Y => \U1/N258\);
    
    \U1/data_all_RNO[97]\ : OA1B
      port map(A => \U1/N_829\, B => \U1/data_filter[1]_net_1\, C
         => \U1/data_all_3_i_0_0_0[97]\, Y => \U1/N_1614\);
    
    \U1/data_all_RNO[88]\ : OA1B
      port map(A => \U1/N_834_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[88]\, Y => \U1/N_202\);
    
    \U2/cnt_RNI767T_0[10]\ : NOR2
      port map(A => \U2/cnt[11]_net_1\, B => \U2/cnt[10]_net_1\, 
        Y => \U2/N_154\);
    
    \U1/data_all_RNO[214]\ : OA1B
      port map(A => \U1/N_840\, B => \U1/data_filter[6]_net_1\, C
         => \U1/data_all_3_0_0_i_0[214]\, Y => \U1/N_182\);
    
    \U2/parity_check_RNO_4\ : OR3
      port map(A => \U2/N_121\, B => \U2/N_119\, C => 
        \U2/parity_check_10_iv_0_1\, Y => 
        \U2/parity_check_10_iv_0_4\);
    
    \U1/data_all_RNO_0[217]\ : NOR2A
      port map(A => \U1/N_840\, B => \data_all[217]\, Y => 
        \U1/N_1019\);
    
    \U5/data_send_RNO_8[4]\ : MX2
      port map(A => \U5/N_375\, B => \U5/N_383\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_479\);
    
    \U5/data_send_RNO_26[2]\ : MX2
      port map(A => \data_all[194]\, B => \data_all[202]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_437\);
    
    \U0/data_ad_RNO[4]\ : NOR2A
      port map(A => \data_in_c[4]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[4]\);
    
    \U5/cnt[3]\ : DFN1E0C0
      port map(D => \U5/cnt_n3\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \U5/cnt[3]_net_1\);
    
    \U1/data_all_RNO_0[234]\ : AO1C
      port map(A => \data_all[234]\, B => \U1/N_837_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[234]\);
    
    \U3/data_recive_RNO_0[2]\ : NOR2A
      port map(A => \data_recive[2]\, B => send_over, Y => 
        \U3/m89_0\);
    
    \U1/pr_state[5]\ : DFN1C0
      port map(D => \U1/N_119\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U1/pr_state[5]_net_1\);
    
    \U2/cnt[1]\ : DFN1C0
      port map(D => \U2/cnt_n1_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[1]_net_1\);
    
    \U5/cnt_RNI6GPF[1]\ : CLKINT
      port map(A => \U5/cnt_0[1]\, Y => \U5/cnt[1]_net_1\);
    
    \U3/un7_cnt_1_I_29\ : AND3
      port map(A => \U3/cnt[6]_net_1\, B => \U3/cnt[7]_net_1\, C
         => \U3/cnt[8]_net_1\, Y => \U3/DWACT_FINC_E[5]\);
    
    \U1/data_all[112]\ : DFN1E0C0
      port map(D => \U1/N_364\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[112]\);
    
    \U3/un7_cnt_1_I_19\ : AND3
      port map(A => \U3/DWACT_FINC_E[0]\, B => 
        \U3/DWACT_FINC_E[2]\, C => \U3/cnt[6]_net_1\, Y => 
        \U3/N_6\);
    
    \U5/data_send_RNO[3]\ : MX2A
      port map(A => \U5/i65_mux\, B => \U5/N_55_0\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[3]\);
    
    \U2/cnt_RNIOPF61[1]\ : OR2
      port map(A => \U2/N_181\, B => \U2/N_180\, Y => 
        \U2/un1_tx_uart27_4_tz\);
    
    \U1/data_all_RNO[137]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[137]\, Y => \U1/N_87\);
    
    \U5/data_send_RNO_25[0]\ : MX2
      port map(A => \data_all[176]\, B => \data_all[184]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_427\);
    
    \U1/m146_i_0_o2_0_0\ : OR2
      port map(A => \U1/m146_i_0_o2_1\, B => \U1/N_817\, Y => 
        \U1/N_838_0\);
    
    \U1/data_all_RNO_0[92]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[92]\, Y => 
        \U1/N_1035\);
    
    \U0/data_ad[6]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[6]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[6]\);
    
    \U1/cnt[2]\ : DFN1E1C0
      port map(D => \U1/cnt_n2_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_793\, Q => \U1/cnt[2]_net_1\);
    
    \U5/data_send_RNO_22[6]\ : MX2
      port map(A => \data_all[134]\, B => \data_all[142]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_409\);
    
    \U3/data_recive[7]\ : DFN1C0
      port map(D => \U3/data_recive_12[7]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[7]\);
    
    \U1/data_all_RNO[228]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_919\, C
         => \U1/N_920\, Y => \U1/N_215\);
    
    \U5/data_send_RNO_27[3]\ : MX2
      port map(A => \data_all[211]\, B => \data_all[219]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_446\);
    
    \U2/cnt_RNIBRJ9[1]\ : NOR2A
      port map(A => \U2/cnt[1]_net_1\, B => \U2/cnt[6]_net_1\, Y
         => \U2/N_163\);
    
    \U1/pr_state_RNO_1[0]\ : NOR2B
      port map(A => \U1/N_854\, B => addr_over, Y => \U1/N_865\);
    
    \U1/data_all_RNO[91]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2131\, C
         => \U1/N_2132\, Y => \U1/N_362\);
    
    \U1/data_all_RNO_1[9]\ : NOR2
      port map(A => \U1/data_filter[9]_net_1\, B => \U1/N_835\, Y
         => \U1/N_1078\);
    
    \U1/data_all_RNO_0[169]\ : AO1C
      port map(A => \data_all[169]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m167_i_0_0\);
    
    \U1/data_all_RNO[197]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m130_0_i_0\, Y => \U1/N_89\);
    
    \U1/data_all[151]\ : DFN1E0C0
      port map(D => \U1/N_130\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[151]\);
    
    \U1/receive_flag\ : DFN1E1C0
      port map(D => addr_over_i, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_263\, Q => \U1/receive_flag_net_1\);
    
    \U1/data_filter_RNO_0[11]\ : AO1D
      port map(A => \U1/data_filter[13]_net_1\, B => 
        \U1/pr_state[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, Y
         => \U1/data_filter_4_i_0_0_0[11]\);
    
    \U1/data_all_RNO_0[166]\ : AO1C
      port map(A => \data_all[166]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m176_i_0_0\);
    
    \U3/cnt_RNIHIT01[6]\ : NOR2B
      port map(A => \U3/N_110_mux\, B => \U3/cnt[6]_net_1\, Y => 
        \U3/N_29\);
    
    \data_in_pad[1]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(1), Y => \data_in_pad[1]/U0/NET1\);
    
    \U1/data_all_RNO_0[162]\ : AO1C
      port map(A => \data_all[162]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m71_i_0_0\);
    
    \U5/data_send[6]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[6]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[6]\);
    
    \U2/cnt_RNI4MI03[10]\ : NOR3C
      port map(A => \U2/N_169\, B => \U2/N_154\, C => 
        \U2/un1_tx_uart27_4_tz\, Y => \U2/un1_tx_uart27_4\);
    
    \U1/data_all_RNO[68]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_971\, C
         => \U1/N_972\, Y => \U1/N_171\);
    
    \U1/data_all[186]\ : DFN1E0C0
      port map(D => \U1/N_413\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[186]\);
    
    \U1/pr_state[1]\ : DFN1C0
      port map(D => \U1/N_867\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U1/pr_state[1]_net_1\);
    
    \U2/send_over\ : DFN1E1C0
      port map(D => \U2/tx_uart38_10\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U2/N_198\, Q => send_over);
    
    \addr_pad[2]/U0/U1\ : IOTRI_OB_EB
      port map(D => \addr_c[2]\, E => \VCC\, DOUT => 
        \addr_pad[2]/U0/NET1\, EOUT => \addr_pad[2]/U0/NET2\);
    
    \U1/data_all_RNO_0[42]\ : NOR2A
      port map(A => \U1/N_832\, B => \data_all[42]\, Y => 
        \U1/N_2199\);
    
    \U1/data_all[174]\ : DFN1E0C0
      port map(D => \U1/data_all_3[174]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[174]\);
    
    \U5/data_send_RNO_4[6]\ : MX2C
      port map(A => \U5/N_497\, B => \U5/N_505\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_531\);
    
    \U1/data_all_RNO_0[168]\ : AO1C
      port map(A => \data_all[168]\, B => \U1/N_838_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m170_i_0_0\);
    
    \U5/data_send_RNO_28[2]\ : MX2
      port map(A => \data_all[226]\, B => \data_all[234]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_453\);
    
    \U5/data_send_RNO_14[3]\ : MX2
      port map(A => \data_all[3]\, B => \data_all[11]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_342\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I70_Y\ : AO1
      port map(A => \U1/N270\, B => \U1/N250\, C => \U1/N269\, Y
         => \U1/N329\);
    
    \U1/cnt_daly_RNO[3]\ : XA1C
      port map(A => \U1/cnt_daly[3]_net_1\, B => \U1/N_846\, C
         => \U1/pr_state[7]_net_1\, Y => \U1/N_800\);
    
    \U0/data_ad_RNO[10]\ : NOR2A
      port map(A => \data_in_c[10]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[10]\);
    
    \U5/data_send[3]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[3]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[3]\);
    
    \U1/data_all_RNO[184]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[184]\, Y => \U1/N_409\);
    
    \U3/un7_cnt_1_I_7\ : AX1C
      port map(A => \U3/cnt[1]_net_1\, B => \U3/cnt[0]_net_1\, C
         => \U3/cnt[2]_net_1\, Y => \U3/I_7\);
    
    \U1/data_all_RNO_0[80]\ : AO1C
      port map(A => \data_all[80]\, B => \U1/N_834_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[80]\);
    
    \U1/data_all[102]\ : DFN1E0C0
      port map(D => \U1/N_54\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[102]\);
    
    \U5/data_send_RNO_9[6]\ : MX2
      port map(A => \U5/N_393\, B => \U5/N_401\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_489\);
    
    \U5/data_send_RNO_3[1]\ : MX2
      port map(A => \U5/N_476\, B => \U5/N_484\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_524\);
    
    \U2/tx_uart_RNO_4\ : AO1
      port map(A => \U2/parity_check_2_sqmuxa\, B => 
        \data_send[1]\, C => \U2/data_send_m[3]\, Y => 
        \U2/tx_uart_11_iv_2\);
    
    \U2/cnt_RNI7NJ9_0[0]\ : NOR2A
      port map(A => \U2/cnt[3]_net_1\, B => \U2/cnt[0]_net_1\, Y
         => \U2/tx_uart35_0_a2_0_0\);
    
    \U1/data_all[49]\ : DFN1E0C0
      port map(D => \U1/N_700\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[49]\);
    
    \U2/idle_send_RNO\ : NOR2A
      port map(A => \U2/send_net_1\, B => \U2/tx_uart38\, Y => 
        \U2/idle_send_0_sqmuxa\);
    
    \U1/data_all[2]\ : DFN1E0C0
      port map(D => \U1/N_2043\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[2]\);
    
    \U1/data_filter_RNO[8]\ : OA1C
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/un2_data_filter[8]\, C => 
        \U1/data_filter_4_i_0_0_0[8]\, Y => \U1/N_39\);
    
    \U1/data_all_RNO_0[121]\ : AO1C
      port map(A => \data_all[121]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[121]\);
    
    \U1/data_all[196]\ : DFN1E0C0
      port map(D => \U1/N_203\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[196]\);
    
    \U1/data_all_RNO[216]\ : OA1B
      port map(A => \U1/N_840_0\, B => \U1/data_filter[8]_net_1\, 
        C => \U1/m64_1_i_0_0\, Y => \U1/N_1779\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I27_Y\ : OA1
      port map(A => \U1/data_filter[5]_net_1\, B => \data_ad[5]\, 
        C => \U1/N189\, Y => \U1/N243\);
    
    \U4/addr_over_RNID0B1\ : INV
      port map(A => addr_over, Y => addr_over_i);
    
    \U5/data_send_RNO_2[4]\ : MX2
      port map(A => \U5/N_463\, B => \U5/N_471\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_519\);
    
    \U1/data_all_RNO[106]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[10]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[106]\, Y => \U1/N_46\);
    
    \U0/cnt_rc[0]\ : DFN1E0C0
      port map(D => \U0/N_164\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/N_135\, Q => \U0/cnt_rc[0]_net_1\);
    
    \U1/data_all_RNO[24]\ : OA1B
      port map(A => \U1/N_836\, B => \U1/data_filter[8]_net_1\, C
         => \U1/m141_0_i_0_0\, Y => \U1/N_1789\);
    
    \addr_pad[1]/U0/U0\ : IOPAD_TRI
      port map(D => \addr_pad[1]/U0/NET1\, E => 
        \addr_pad[1]/U0/NET2\, PAD => addr(1));
    
    \U0/data_ad_RNO[1]\ : NOR2A
      port map(A => \data_in_c[1]\, B => \U0/pr_state[5]_net_1\, 
        Y => \U0/data_ad_4[1]\);
    
    \U3/cnt_RNI3VAQ1[2]\ : NOR3C
      port map(A => \U3/m17_1\, B => \U3/m17_0\, C => 
        \U3/N_110_mux\, Y => \U3/N_125_mux\);
    
    \U5/data_send_RNO_7[7]\ : MX2
      port map(A => \U5/N_362\, B => \U5/N_370\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_474\);
    
    \U1/data_all[189]\ : DFN1E0C0
      port map(D => \U1/N_419\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[189]\);
    
    \U5/data_send_RNO_17[4]\ : MX2
      port map(A => \data_all[52]\, B => \data_all[60]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_367\);
    
    \U2/cnt_c2\ : NOR3C
      port map(A => \U2/cnt[1]_net_1\, B => \U2/cnt[0]_net_1\, C
         => \U2/cnt[2]_net_1\, Y => \U2/cnt_c2_net_1\);
    
    \U2/cnt_RNI7DUF2_0[1]\ : NOR2B
      port map(A => \U2/N_196\, B => \U2/N_173\, Y => 
        \U2/parity_check_2_sqmuxa\);
    
    \U4/addr_RNO[2]\ : XA1
      port map(A => \addr_c[2]\, B => \U4/N_8_0\, C => 
        \U4/pr_state[0]_net_1\, Y => \U4/addr_n2\);
    
    \U3/data_recive_RNO[2]\ : MX2
      port map(A => \U3/m89_0\, B => rx_uart_c, S => 
        \U3/data_recive25\, Y => \U3/data_recive_12[2]\);
    
    \U1/data_all_RNO_1[145]\ : NOR2
      port map(A => \U1/data_filter[1]_net_1\, B => \U1/N_842\, Y
         => \U1/N_2248\);
    
    \U1/data_all_RNO[17]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2275\, C
         => \U1/N_2276\, Y => \U1/N_1783\);
    
    \U1/data_all_RNO_0[210]\ : AO1C
      port map(A => \data_all[210]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[210]\);
    
    \U4/addr[1]\ : DFN1E0C0
      port map(D => \U4/addr_n1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U4/N_7_0\, Q => \addr_c[1]\);
    
    \U1/data_filter_RNO_0[7]\ : AO1D
      port map(A => \U1/data_filter[9]_net_1\, B => 
        \U1/pr_state[5]_net_1\, C => \U1/pr_state[7]_net_1\, Y
         => \U1/m48_0_0_0\);
    
    \U1/data_filter[3]\ : DFN1E0C0
      port map(D => \U1/N_1421\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[3]_net_1\);
    
    \U1/data_all_RNO_0[71]\ : AO1C
      port map(A => \data_all[71]\, B => \U1/N_833\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m231_i_0_0\);
    
    \U1/data_filter[4]\ : DFN1E0C0
      port map(D => \U1/N_41\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[4]_net_1\);
    
    \U1/data_all_RNO[202]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_925\, C
         => \U1/N_926\, Y => \U1/N_77\);
    
    \U1/cnt_daly_RNO[9]\ : XA1B
      port map(A => \U1/m24_N_11_mux\, B => 
        \U1/cnt_daly[9]_net_1\, C => \U1/pr_state_0[7]_net_1\, Y
         => \U1/cnt_daly_n9\);
    
    \U4/addr_RNI62K31[0]\ : OA1C
      port map(A => \U4.N_31\, B => \addr_c[0]\, C => 
        ad_once_over, Y => \U4/N_6_0\);
    
    \U1/data_all_RNO_0[208]\ : AO1C
      port map(A => \data_all[208]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[208]\);
    
    \U1/pr_state_RNICDI39[1]\ : OR3
      port map(A => \U1/N_866\, B => \U1/pr_state[1]_net_1\, C
         => \U1/N_871\, Y => \U1/pr_state_RNICDI39[1]_net_1\);
    
    \U1/data_all_RNO[73]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[9]_net_1\, 
        C => \U1/m225_i_0_0\, Y => \U1/N_181\);
    
    \U5/data_send_RNO_9[3]\ : MX2
      port map(A => \U5/N_390\, B => \U5/N_398\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_486\);
    
    \U2/cnt_RNISS7J_0[1]\ : NOR3A
      port map(A => \U2/un1_tx_uart27_3_0_a2_3_0\, B => 
        \U2/cnt[6]_net_1\, C => \U2/cnt[1]_net_1\, Y => 
        \U2/un1_tx_uart27_3_0_a2_3_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I80_Y\ : AO1
      port map(A => \U1/N271\, B => \U1/N264\, C => 
        \U1/ADD_14x14_fast_I80_Y_0\, Y => \U1/N321\);
    
    \U1/pr_state[4]\ : DFN1C0
      port map(D => \U1/pr_state_ns[3]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U1/pr_state[4]_net_1\);
    
    \sts_pad/U0/U1\ : IOIN_IB
      port map(YIN => \sts_pad/U0/NET1\, Y => sts_c);
    
    \U1/data_all_RNO_0[184]\ : AO1C
      port map(A => \data_all[184]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[184]\);
    
    \U1/data_all_RNO_0[173]\ : AO1C
      port map(A => \data_all[173]\, B => \U1/N_838_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m153_i_0_0\);
    
    \data_in_pad[2]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(2), Y => \data_in_pad[2]/U0/NET1\);
    
    \U5/data_send_RNO_24[4]\ : MX2
      port map(A => \data_all[164]\, B => \data_all[172]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_423\);
    
    \U5/data_send_RNO_15[7]\ : MX2
      port map(A => \data_all[23]\, B => \data_all[31]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_354\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I23_Y\ : OA1
      port map(A => \U1/data_filter[7]_net_1\, B => \data_ad[7]\, 
        C => \U1/N195\, Y => \U1/N239\);
    
    \U3/data_recive_RNO_3[6]\ : NOR3B
      port map(A => \U3/cnt[10]_net_1\, B => \U3/cnt[3]_net_1\, C
         => \U3/cnt[7]_net_1\, Y => \U3/m79_3\);
    
    \U1/data_all_RNO[103]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[7]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[103]\, Y => \U1/N_52\);
    
    \U5/data_send_RNO_26[3]\ : MX2
      port map(A => \data_all[195]\, B => \data_all[203]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_438\);
    
    \U1/cnt_daly_RNITBVQ[4]\ : NOR2B
      port map(A => \U1/cnt_daly[4]_net_1\, B => 
        \U1/cnt_daly[5]_net_1\, Y => \U1/m20_m6_0_a2_2\);
    
    \U2/tx_uart_RNO\ : OR3
      port map(A => \U2/tx_uart_11_iv_6\, B => 
        \U2/tx_uart_11_iv_5\, C => \U2/tx_uart_11_iv_7\, Y => 
        \U2/tx_uart_11\);
    
    \U2/cnt_RNIULDJ[9]\ : NOR2
      port map(A => \U2/cnt[9]_net_1\, B => \U2/cnt[10]_net_1\, Y
         => \U2/tx_uart37_6\);
    
    \U2/cnt_RNI8PAD2_0[1]\ : NOR3C
      port map(A => \U2/N_171\, B => 
        \U2/un1_tx_uart27_3_0_a2_3_1\, C => \U2/tx_uart34_1\, Y
         => \U2/N_111\);
    
    \U1/data_all[199]\ : DFN1E0C0
      port map(D => \U1/N_85\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[199]\);
    
    \U5/data_send_RNO[0]\ : MX2A
      port map(A => \U5/i59_mux\, B => \U5/N_76\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[0]\);
    
    \U2/cnt_RNIH1K9[8]\ : NOR2B
      port map(A => \U2/cnt[8]_net_1\, B => \U2/cnt[5]_net_1\, Y
         => \U2/N_129\);
    
    \U1/data_all_RNO_0[177]\ : AO1C
      port map(A => \data_all[177]\, B => \U1/N_844_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[177]\);
    
    \U1/data_all_RNO[100]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[100]\, Y => \U1/N_58\);
    
    \U1/delay_channel1_RNO_1\ : NOR2A
      port map(A => \U1/pr_state[1]_net_1\, B => 
        \U1/pr_state[0]_net_1\, Y => \U1/N_872\);
    
    \U1/data_all_RNO[112]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[112]\, Y => \U1/N_364\);
    
    \U1/data_all_RNO[4]\ : OA1B
      port map(A => \U1/N_835_0\, B => \U1/data_filter[4]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[4]\, Y => \U1/N_255\);
    
    \U1/data_all_RNO[11]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1075\, C
         => \U1/N_1076\, Y => \U1/N_241\);
    
    \U1/data_all[111]\ : DFN1E0C0
      port map(D => \U1/N_1608\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[111]\);
    
    \addr_pad[0]/U0/U0\ : IOPAD_TRI
      port map(D => \addr_pad[0]/U0/NET1\, E => 
        \addr_pad[0]/U0/NET2\, PAD => addr(0));
    
    \U1/data_filter_RNO_0[9]\ : AO1D
      port map(A => \U1/data_filter[11]_net_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, 
        Y => \U1/m45_0_0_0\);
    
    \U5/data_send_RNO_7[1]\ : MX2
      port map(A => \U5/N_356\, B => \U5/N_364\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_468\);
    
    \U1/data_all_RNO[239]\ : NOR3C
      port map(A => \data_all[239]\, B => \U1/pr_state[2]_net_1\, 
        C => \U1/N_837\, Y => \U1/N_252\);
    
    \U1/m302_0_i_o2_0\ : OR3A
      port map(A => \addr_c_0[0]\, B => \U1/I_5_0\, C => 
        \U1/I_9_0\, Y => \U1/m302_0_i_o2_0_net_1\);
    
    \U1/data_all_RNO_0[36]\ : AO1C
      port map(A => \data_all[36]\, B => \U1/N_832_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m286_i_0_0\);
    
    \U5/data_send_RNO_12[0]\ : MX2
      port map(A => \U5/N_435\, B => \U5/N_443\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_507\);
    
    \U5/data_send_RNO[5]\ : MX2A
      port map(A => \U5/i69_mux\, B => \U5/N_41_0\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[5]\);
    
    \U1/data_all[158]\ : DFN1E0C0
      port map(D => \U1/data_all_3[158]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[158]\);
    
    \U1/receive_on_RNO\ : AO1
      port map(A => \U1/m110_i_0_a3_1\, B => \U1/N_139\, C => 
        addr_over, Y => \U1/N_260\);
    
    \U1/data_all_RNO_0[147]\ : AO1C
      port map(A => \data_all[147]\, B => \U1/N_842_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m109_0_i_0_0\);
    
    \U1/data_all_RNO[83]\ : OA1B
      port map(A => \U1/N_834_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[83]\, Y => \U1/N_212\);
    
    \U0/sts_ris3\ : DFN1C0
      port map(D => \U0/sts_ris2_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U0/sts_ris3_net_1\);
    
    \U3/data_recive_RNO_4[6]\ : NOR2B
      port map(A => \U3/cnt[1]_net_1\, B => \U3/cnt[0]_net_1\, Y
         => \U3/m79_2\);
    
    \U1/data_all_RNO_0[39]\ : NOR2A
      port map(A => \U1/N_832\, B => \data_all[39]\, Y => 
        \U1/N_2205\);
    
    \U5/data_send_RNO_6[7]\ : MX2
      port map(A => \U5/N_346\, B => \U5/N_354\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_466\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I4_P0N\ : OR2
      port map(A => \data_ad[4]\, B => \U1/data_filter[4]_net_1\, 
        Y => \U1/N189\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I18_Y\ : AO1
      port map(A => \U1/N200\, B => \U1/N204\, C => \U1/N203\, Y
         => \U1/N234\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I15_Y\ : OA1
      port map(A => \U1/data_filter[11]_net_1\, B => 
        \data_ad[11]\, C => \U1/N207\, Y => \U1/N231\);
    
    \U1/data_all_RNO_0[204]\ : AO1C
      port map(A => \data_all[204]\, B => \U1/N_839_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[204]\);
    
    \U2/cnt_c1_i\ : OR2B
      port map(A => \U2/cnt[0]_net_1\, B => \U2/cnt[1]_net_1\, Y
         => \U2/N_7\);
    
    \U5/data_send_RNO_17[6]\ : MX2
      port map(A => \data_all[54]\, B => \data_all[62]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_369\);
    
    \U4/addr[3]\ : DFN1E0C0
      port map(D => \U4/addr_n3\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U4/N_7_0\, Q => \addr_c[3]\);
    
    \U3/cnt_4[7]\ : XA1
      port map(A => \U3/N_6\, B => \U3/cnt[7]_net_1\, C => 
        \U3/recive_net_1\, Y => \U3/cnt_4[7]_net_1\);
    
    \U1/cnt_daly_RNO_3[10]\ : NOR2B
      port map(A => \U1/cnt_daly[5]_net_1\, B => 
        \U1/cnt_daly[6]_net_1\, Y => \U1/m22_m4_0_a2_2\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I10_G0N\ : NOR2B
      port map(A => \data_ad[10]\, B => 
        \U1/data_filter[10]_net_1\, Y => \U1/N206\);
    
    \U5/data_send_RNO_1[1]\ : MX2A
      port map(A => \U5/N_536\, B => \U5/N_68\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_69\);
    
    \U1/data_filter_RNO[1]\ : OA1C
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/un2_data_filter[1]\, C => \U1/m57_0_0_0\, Y => 
        \U1/N_58_0\);
    
    \U1/data_all[217]\ : DFN1E0C0
      port map(D => \U1/N_174\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[217]\);
    
    \rc_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => rc_c, E => \VCC\, DOUT => \rc_pad/U0/NET1\, 
        EOUT => \rc_pad/U0/NET2\);
    
    \U5/data_send_RNO_17[7]\ : MX2
      port map(A => \data_all[55]\, B => \data_all[63]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_370\);
    
    \U1/data_all_RNO[134]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[134]\, Y => \U1/N_82\);
    
    \U0/conver_ris3_RNO\ : INV
      port map(A => \U0/conver_ris2_net_1\, Y => 
        \U0/conver_ris2_i\);
    
    \U5/data_send_RNO_9[1]\ : MX2
      port map(A => \U5/N_388\, B => \U5/N_396\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_484\);
    
    \U5/data_send_RNO_28[5]\ : MX2
      port map(A => \data_all[229]\, B => \data_all[237]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_456\);
    
    \U1/data_all_RNO[231]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_985\, C
         => \U1/N_986\, Y => \U1/N_32\);
    
    \U1/data_all_RNO_0[160]\ : AO1C
      port map(A => \data_all[160]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m191_i_0_0\);
    
    \U1/data_all[73]\ : DFN1E0C0
      port map(D => \U1/N_181\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[73]\);
    
    \U1/cnt_daly_RNO_2[9]\ : NOR3C
      port map(A => \U1/cnt_daly[5]_net_1\, B => 
        \U1/cnt_daly[2]_net_1\, C => \U1/cnt_daly[7]_net_1\, Y
         => \U1/m24_m4_e_3\);
    
    \U1/data_all_RNO[142]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[142]\, 
        C => \U1/N_841_0\, Y => \U1/N_19\);
    
    \U3/cnt_RNIFBUG[8]\ : NOR2A
      port map(A => \U3/cnt[1]_net_1\, B => \U3/cnt[8]_net_1\, Y
         => \U3/m27_1\);
    
    \U2/cnt_RNI6QQV[10]\ : NOR3B
      port map(A => \U2/send_net_1\, B => \U2/cnt[10]_net_1\, C
         => \U2/cnt[11]_net_1\, Y => \U2/N_168\);
    
    \U1/data_all_RNO_0[96]\ : AO1C
      port map(A => \data_all[96]\, B => \U1/N_829_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[96]\);
    
    \U1/data_all_RNO_0[99]\ : AO1C
      port map(A => \data_all[99]\, B => \U1/N_829_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[99]\);
    
    \U1/data_filter[1]\ : DFN1E0C0
      port map(D => \U1/N_58_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[1]_net_1\);
    
    \U1/data_all_RNO[90]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2291\, C
         => \U1/N_2292\, Y => \U1/N_1775\);
    
    \U1/data_all_RNO[230]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_915\, C
         => \U1/N_916\, Y => \U1/N_219\);
    
    \U1/data_all_RNO[129]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[1]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[129]\, Y => \U1/N_73\);
    
    \U5/data_send_RNO_13[1]\ : NOR2A
      port map(A => \U5/N_452\, B => \U5/cnt[1]_net_1\, Y => 
        \U5/N_67_0\);
    
    \U1/m125_0_0_i_o2_0\ : OR3
      port map(A => \addr_c_0[0]\, B => \U1/I_5_0\, C => 
        \U1/I_9_0\, Y => \U1/m125_0_0_i_o2_0_net_1\);
    
    \U1/data_all_RNO[194]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/m139_0_i_0\, Y => \U1/N_93\);
    
    \U0/pr_state[5]\ : DFN1P0
      port map(D => \U0/pr_state_ns[0]\, CLK => sys_clk_c, PRE
         => sys_rest_c, Q => \U0/pr_state[5]_net_1\);
    
    \data_in_pad[6]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(6), Y => \data_in_pad[6]/U0/NET1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I51_Y\ : NOR2B
      port map(A => \U1/N247\, B => \U1/N243\, Y => \U1/N270\);
    
    \U1/data_all_RNO_0[83]\ : AO1C
      port map(A => \data_all[83]\, B => \U1/N_834_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[83]\);
    
    \U1/data_all[136]\ : DFN1E0C0
      port map(D => \U1/N_103\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[136]\);
    
    \U1/data_all_RNO_0[115]\ : AO1C
      port map(A => \data_all[115]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[115]\);
    
    \cs_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \GND\, E => \VCC\, DOUT => \cs_pad/U0/NET1\, 
        EOUT => \cs_pad/U0/NET2\);
    
    \U5/data_send_RNO_0[4]\ : MX2C
      port map(A => \U5/N_519\, B => \U5/N_527\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i67_mux\);
    
    \U1/data_all_RNO[63]\ : NOR3C
      port map(A => \data_all[63]\, B => \U1/pr_state[2]_net_1\, 
        C => \U1/N_831\, Y => \U1/N_91\);
    
    \U1/un14_data_all_I_8\ : OR3
      port map(A => \addr_c_0[0]\, B => \addr_c[1]\, C => 
        \addr_c[2]\, Y => \U1/N_3\);
    
    \U1/data_all[101]\ : DFN1E0C0
      port map(D => \U1/N_56\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[101]\);
    
    \U5/data_send_RNO_22[1]\ : MX2
      port map(A => \data_all[129]\, B => \data_all[137]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_404\);
    
    \U1/data_all_RNO_1[228]\ : NOR2
      port map(A => \U1/data_filter[4]_net_1\, B => \U1/N_837\, Y
         => \U1/N_920\);
    
    \U1/data_all_RNO_0[52]\ : AO1C
      port map(A => \data_all[52]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[52]\);
    
    \U1/data_all_RNO[72]\ : OA1B
      port map(A => \U1/N_833\, B => \U1/data_filter[8]_net_1\, C
         => \U1/m228_i_0_0\, Y => \U1/N_179\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I43_Y\ : NOR2B
      port map(A => \U1/N239\, B => \U1/N235\, Y => \U1/N262\);
    
    \U5/data_send_RNO_23[6]\ : MX2
      port map(A => \data_all[150]\, B => \data_all[158]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_417\);
    
    \U1/data_all_RNO[208]\ : OA1B
      port map(A => \U1/N_840_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[208]\, Y => \U1/N_196\);
    
    \U5/data_send_RNO_1[3]\ : MX2A
      port map(A => \U5/N_534\, B => \U5/N_54_0\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_55_0\);
    
    \U1/data_all_RNO[188]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[188]\, Y => \U1/N_417\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I79_un1_Y\ : NOR3C
      port map(A => \U1/N270\, B => \U1/N262\, C => \U1/N250\, Y
         => \U1/I79_un1_Y\);
    
    \U1/data_all_RNO_0[49]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[49]\, Y => 
        \U1/N_2155\);
    
    \U5/data_send_RNO_11[6]\ : MX2
      port map(A => \U5/N_425\, B => \U5/N_433\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_505\);
    
    \U1/cnt_daly_RNO[4]\ : NOR3A
      port map(A => \U1/N_848\, B => \U1/N_2299\, C => 
        \U1/pr_state[7]_net_1\, Y => \U1/N_802\);
    
    \U1/data_all[207]\ : DFN1E0C0
      port map(D => \U1/N_158\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[207]\);
    
    \U1/data_all[145]\ : DFN1E0C0
      port map(D => \U1/N_1795\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[145]\);
    
    \U5/data_send_RNO_19[6]\ : MX2
      port map(A => \data_all[86]\, B => \data_all[94]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_385\);
    
    \U5/data_send_RNO_16[0]\ : MX2
      port map(A => \data_all[32]\, B => \data_all[40]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_355\);
    
    \U1/cnt_daly_RNO[1]\ : XA1B
      port map(A => \U1/cnt_daly[0]_net_1\, B => 
        \U1/cnt_daly[1]_net_1\, C => \U1/pr_state_0[7]_net_1\, Y
         => \U1/N_796\);
    
    \U5/data_send_RNO_25[4]\ : MX2
      port map(A => \data_all[180]\, B => \data_all[188]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_431\);
    
    \U5/data_send_RNO_24[5]\ : MX2
      port map(A => \data_all[165]\, B => \data_all[173]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_424\);
    
    \U2/cnt[0]\ : DFN1C0
      port map(D => \U2/cnt_n0_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[0]_net_1\);
    
    \U0/pr_state[1]\ : DFN1C0
      port map(D => \U0/pr_state[2]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U0/pr_state[1]_net_1\);
    
    \U5/data_send_RNO_22[4]\ : MX2
      port map(A => \data_all[132]\, B => \data_all[140]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_407\);
    
    \U1/data_all_RNO_0[67]\ : AO1C
      port map(A => \data_all[67]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m243_i_0_0\);
    
    \U1/data_all_RNO[82]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1047\, C
         => \U1/N_1048\, Y => \U1/N_216\);
    
    \U1/data_all[165]\ : DFN1E0C0
      port map(D => \U1/N_317\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[165]\);
    
    \U2/cnt_RNI919L1[9]\ : NOR3C
      port map(A => \U2/un1_cnt_2\, B => \U2/un1_cnt_1\, C => 
        \U2/un1_cnt_5\, Y => \U2/un1_cnt_8\);
    
    \U5/data_send_RNO_21[5]\ : MX2
      port map(A => \data_all[117]\, B => \data_all[125]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_400\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I6_G0N\ : NOR2B
      port map(A => \data_ad[6]\, B => \U1/data_filter[6]_net_1\, 
        Y => \U1/N194\);
    
    \U1/data_filter_RNO[6]\ : OA1C
      port map(A => \U1/pr_state_0[5]_net_1\, B => 
        \U1/un2_data_filter[6]\, C => \U1/m51_0_0_0\, Y => 
        \U1/N_52_0\);
    
    \U3/cnt[3]\ : DFN1C0
      port map(D => \U3/cnt_4[3]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U3/cnt[3]_net_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I6_P0N\ : OR2
      port map(A => \data_ad[6]\, B => \U1/data_filter[6]_net_1\, 
        Y => \U1/N195\);
    
    \U1/data_all_3_i_o2_i_a3_i_o2_0_o2[63]\ : OR2
      port map(A => 
        \U1/data_all_3_i_o2_i_a3_i_o2_0_o2_0[63]_net_1\, B => 
        \U1/N_817\, Y => \U1/N_831\);
    
    \U1/data_all[212]\ : DFN1E0C0
      port map(D => \U1/N_190\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[212]\);
    
    \U5/data_send_RNO_9[2]\ : MX2
      port map(A => \U5/N_389\, B => \U5/N_397\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_485\);
    
    \U1/data_all[126]\ : DFN1E0C0
      port map(D => \U1/N_72\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[126]\);
    
    \U1/data_all_RNO_0[119]\ : AO1C
      port map(A => \data_all[119]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[119]\);
    
    \U1/data_all[239]\ : DFN1E0C0
      port map(D => \U1/N_252\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[239]\);
    
    \U5/data_send_RNO_28[7]\ : MX2
      port map(A => \data_all[231]\, B => \data_all[239]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_458\);
    
    \U1/data_all_RNO_0[27]\ : NOR2A
      port map(A => \U1/N_836\, B => \data_all[27]\, Y => 
        \U1/N_2255\);
    
    \U1/data_all_RNO_0[116]\ : AO1C
      port map(A => \data_all[116]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[116]\);
    
    \U3/cnt[7]\ : DFN1C0
      port map(D => \U3/cnt_4[7]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U3/cnt[7]_net_1\);
    
    \U1/data_all[78]\ : DFN1E0C0
      port map(D => \U1/data_all_3[78]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[78]\);
    
    \U1/data_all_RNO_0[112]\ : AO1C
      port map(A => \data_all[112]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[112]\);
    
    \U1/data_all_RNO_0[84]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[84]\, Y => 
        \U1/N_1043\);
    
    \U1/data_all[139]\ : DFN1E0C0
      port map(D => \U1/N_1837\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[139]\);
    
    \U1/data_all[154]\ : DFN1E0C0
      port map(D => \U1/N_1800\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[154]\);
    
    \U1/data_all_RNO[34]\ : OA1B
      port map(A => \U1/N_832\, B => \U1/data_filter[2]_net_1\, C
         => \U1/m292_i_0_0\, Y => \U1/N_1807\);
    
    \U1/cnt_daly[5]\ : DFN1E0C0
      port map(D => \U1/N_804\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[5]_net_1\);
    
    \U1/pr_state[0]\ : DFN1C0
      port map(D => \U1/pr_state_RNO[0]_net_1\, CLK => sys_clk_c, 
        CLR => sys_rest_c, Q => \U1/pr_state[0]_net_1\);
    
    \U1/data_all_RNO_0[118]\ : AO1C
      port map(A => \data_all[118]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[118]\);
    
    \U4/nx_state_RNO[1]\ : MX2A
      port map(A => \U4/N_24\, B => \U4/N_25\, S => 
        \U4/pr_state[0]_net_1\, Y => \U4/nx_state_RNO[1]_net_1\);
    
    \U1/data_all_RNO[115]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[115]\, Y => \U1/N_370\);
    
    \U1/data_all[118]\ : DFN1E0C0
      port map(D => \U1/N_376\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[118]\);
    
    \U1/cnt_daly_RNIVMPM1[1]\ : NOR3A
      port map(A => \U1/m61_0_i_a3_1_2\, B => 
        \U1/cnt_daly[0]_net_1\, C => \U1/cnt_daly[1]_net_1\, Y
         => \U1/m61_0_i_a3_1_7\);
    
    \U1/pr_state_RNIS9HE[3]\ : NOR2A
      port map(A => \U1/pr_state[3]_net_1\, B => send_whole_over, 
        Y => \U1/N_858\);
    
    \U1/data_filter_RNO_0[10]\ : AO1D
      port map(A => \U1/data_filter[12]_net_1\, B => 
        \U1/pr_state[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, Y
         => \U1/data_filter_4_i_0_0_0[10]\);
    
    \U1/data_all_RNO_0[65]\ : AO1C
      port map(A => \data_all[65]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m249_i_0_0\);
    
    \U1/data_all_RNO[62]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[62]\, 
        C => \U1/N_831_0\, Y => \U1/N_1422\);
    
    \U4/addr_RNILUJF[1]\ : NOR2B
      port map(A => \addr_c[1]\, B => \addr_c[0]\, Y => 
        \U4/N_8_0\);
    
    \U1/data_all_RNO_0[70]\ : AO1C
      port map(A => \data_all[70]\, B => \U1/N_833_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m234_i_0_0\);
    
    \U5/data_send_RNO_28[3]\ : MX2
      port map(A => \data_all[227]\, B => \data_all[235]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_454\);
    
    \U5/cnt[4]\ : DFN1E0C0
      port map(D => \U5/cnt_n4\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \U5/cnt[4]_net_1\);
    
    \U2/cnt_n10\ : XA1
      port map(A => \U2/cnt_c9_net_1\, B => \U2/cnt[10]_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n10_net_1\);
    
    \U3/data_recive_RNO_1[6]\ : NOR3C
      port map(A => \U3/m79_4\, B => \U3/m79_3\, C => \U3/N_30_0\, 
        Y => \U3/data_recive29\);
    
    \U1/pr_state_RNO[3]\ : OA1B
      port map(A => \U1/N_857\, B => \U1/N_858\, C => 
        \U1/m68_i_i_1\, Y => \U1/pr_state_RNO[3]_net_1\);
    
    \U1/data_all_RNO_0[4]\ : AO1C
      port map(A => \data_all[4]\, B => \U1/N_835_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[4]\);
    
    \U1/pr_state_RNO[1]\ : NOR2B
      port map(A => send_whole_over, B => \U1/pr_state[3]_net_1\, 
        Y => \U1/N_867\);
    
    \U1/m206_i_0_o2_0_0\ : OR2
      port map(A => \U1/N_826\, B => \U1/N_819\, Y => 
        \U1/N_833_0\);
    
    \U5/data_send_RNO_10[3]\ : MX2
      port map(A => \U5/N_406\, B => \U5/N_414\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_494\);
    
    \U2/cnt_RNIPGDJ[10]\ : NOR2A
      port map(A => \U2/cnt[4]_net_1\, B => \U2/cnt[10]_net_1\, Y
         => \U2/un1_cnt_2\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I21_Y\ : OA1
      port map(A => \U1/data_filter[7]_net_1\, B => \data_ad[7]\, 
        C => \U1/N201\, Y => \U1/N237\);
    
    \U1/data_all_RNO_0[5]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[5]\, Y => 
        \U1/N_1086\);
    
    \U1/data_all[229]\ : DFN1E0C0
      port map(D => \U1/N_217\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[229]\);
    
    \U1/data_all[72]\ : DFN1E0C0
      port map(D => \U1/N_179\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[72]\);
    
    \U1/data_all_RNO_0[25]\ : AO1C
      port map(A => \data_all[25]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m138_0_i_0_0\);
    
    \U1/pr_state_RNIV2MS_0[1]\ : CLKINT
      port map(A => \U1/pr_state_RNIV2MS[1]_net_1\, Y => 
        \U1/N_1091\);
    
    \U1/data_all[202]\ : DFN1E0C0
      port map(D => \U1/N_77\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[202]\);
    
    \U2/cnt_RNIOO7J_0[8]\ : NOR2B
      port map(A => \U2/N_129\, B => \U2/N_165\, Y => \U2/N_153\);
    
    \U5/data_send_RNO_27[0]\ : MX2
      port map(A => \data_all[208]\, B => \data_all[216]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_443\);
    
    \U2/cnt_RNIUU7J[2]\ : NOR3A
      port map(A => \U2/N_176\, B => \U2/cnt[2]_net_1\, C => 
        \U2/cnt[7]_net_1\, Y => \U2/tx_uart27_0_a2_1\);
    
    \U1/data_all[129]\ : DFN1E0C0
      port map(D => \U1/N_73\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[129]\);
    
    \U1/data_all_RNO_0[181]\ : AO1C
      port map(A => \data_all[181]\, B => \U1/N_844\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[181]\);
    
    \U1/data_all_RNO[145]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2247\, C
         => \U1/N_2248\, Y => \U1/N_1795\);
    
    \U1/data_all_RNO[10]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2295\, C
         => \U1/N_2296\, Y => \U1/N_789\);
    
    \U1/data_all_RNO[75]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_957\, C
         => \U1/N_958\, Y => \U1/N_185\);
    
    \U1/m125_0_0_i_o2_0_0\ : OR2
      port map(A => \U1/m125_0_0_i_o2_0_net_1\, B => \U1/N_817\, 
        Y => \U1/N_836_0\);
    
    \U2/cnt_0_sqmuxa\ : NOR2A
      port map(A => \U2/send_net_1\, B => \U2/un1_cnt\, Y => 
        \U2/cnt_0_sqmuxa_net_1\);
    
    \U5/data_send_RNO_4[5]\ : MX2C
      port map(A => \U5/N_496\, B => \U5/N_504\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_116\);
    
    \U1/data_all_RNO_0[219]\ : NOR2A
      port map(A => \U1/N_840\, B => \data_all[219]\, Y => 
        \U1/N_1017\);
    
    \U1/cnt_daly_RNIAJQR[2]\ : NOR2A
      port map(A => \U1/pr_state[0]_net_1\, B => 
        \U1/cnt_daly[2]_net_1\, Y => \U1/m61_0_i_a3_1_2\);
    
    \U0/pr_state[4]\ : DFN1C0
      port map(D => \U0/pr_state_ns[1]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U0/pr_state[4]_net_1\);
    
    \U1/data_all_RNO[235]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_909\, C
         => \U1/N_910\, Y => \U1/N_225\);
    
    \U5/send_whole_over_RNO\ : MX2A
      port map(A => \U5/pr_state[0]_net_1\, B => \U5/N_138_mux\, 
        S => \U5/pr_state[1]_net_1\, Y => \U5/un1_pr_state_1\);
    
    \U3/data_recive_RNO_3[0]\ : NOR3B
      port map(A => \U3/cnt[0]_net_1\, B => \U3/m62_4\, C => 
        \U3/cnt[1]_net_1\, Y => \U3/m62_6\);
    
    \U1/data_all_RNO_1[138]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_841\, 
        Y => \U1/N_948\);
    
    \U1/data_all[108]\ : DFN1E0C0
      port map(D => \U1/N_1611\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[108]\);
    
    \U5/data_send_RNO_10[1]\ : MX2
      port map(A => \U5/N_404\, B => \U5/N_412\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_492\);
    
    \U1/data_all_RNO[138]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_947\, C
         => \U1/N_948\, Y => \U1/N_101\);
    
    \U1/data_all_RNO[181]\ : OA1B
      port map(A => \U1/N_844_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[181]\, Y => \U1/N_403\);
    
    \U3/data_recive[4]\ : DFN1C0
      port map(D => \U3/data_recive_12[4]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[4]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I96_Y_0\ : XOR2
      port map(A => \data_ad[8]\, B => \U1/data_filter[8]_net_1\, 
        Y => \U1/ADD_14x14_fast_I96_Y_0\);
    
    \U3/receive_over_RNO\ : NOR2A
      port map(A => \U3/recive_net_1\, B => \U3/data_recive31\, Y
         => \U3/receive_over_0_sqmuxa\);
    
    \U1/data_all_RNO[85]\ : OA1B
      port map(A => \U1/N_834_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[85]\, Y => \U1/N_208\);
    
    \U1/data_all[71]\ : DFN1E0C0
      port map(D => \U1/N_177\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[71]\);
    
    \U5/data_send_RNO_0[1]\ : MX2C
      port map(A => \U5/N_516\, B => \U5/N_524\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i61_mux\);
    
    \U1/data_all_RNO_0[228]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[228]\, Y => 
        \U1/N_919\);
    
    \U1/data_all_RNO_1[84]\ : NOR2
      port map(A => \U1/data_filter[4]_net_1\, B => \U1/N_834\, Y
         => \U1/N_1044\);
    
    \U1/data_all_RNO_1[231]\ : NOR2
      port map(A => \U1/data_filter[7]_net_1\, B => \U1/N_837\, Y
         => \U1/N_986\);
    
    \U1/data_all[77]\ : DFN1E0C0
      port map(D => \U1/N_724\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[77]\);
    
    \data_in_pad[3]/U0/U0\ : IOPAD_IN
      port map(PAD => data_in(3), Y => \data_in_pad[3]/U0/NET1\);
    
    \U5/data_send_RNO_11[4]\ : MX2
      port map(A => \U5/N_423\, B => \U5/N_431\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_503\);
    
    \U1/data_filter[13]\ : DFN1E0C0
      port map(D => \U1/data_filter_4[13]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[13]_net_1\);
    
    \U1/data_all_RNO[117]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[117]\, Y => \U1/N_374\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I9_G0N\ : NOR2B
      port map(A => \data_ad[9]\, B => \U1/data_filter[9]_net_1\, 
        Y => \U1/N203\);
    
    \U1/data_all_RNO_1[11]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_835\, 
        Y => \U1/N_1076\);
    
    \U1/data_all_RNO[198]\ : OA1B
      port map(A => \U1/N_839_0\, B => \U1/data_filter[6]_net_1\, 
        C => \U1/m127_i_0_0\, Y => \U1/N_206\);
    
    \U1/data_filter_RNO_0[5]\ : AO1D
      port map(A => \U1/data_filter[7]_net_1\, B => 
        \U1/pr_state[5]_net_1\, C => \U1/pr_state[7]_net_1\, Y
         => \U1/m54_0_0_0\);
    
    \U1/cnt_daly_RNIREDU2[6]\ : OR2A
      port map(A => \U1/cnt_daly[6]_net_1\, B => \U1/N_849\, Y
         => \U1/N_850\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I1_P0N\ : OR2
      port map(A => \data_ad[1]\, B => \U1/data_filter[1]_net_1\, 
        Y => \U1/N180\);
    
    \U5/data_send_RNO_0[3]\ : MX2C
      port map(A => \U5/N_518\, B => \U5/N_526\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i65_mux\);
    
    \U3/data_recive_RNO_1[5]\ : NOR3C
      port map(A => \U3/m47_3\, B => \U3/m47_2\, C => 
        \U3/N_120_mux\, Y => \U3/data_recive28\);
    
    \U1/pr_state_RNO_1[6]\ : NOR3A
      port map(A => \U1/pr_state[6]_net_1\, B => ad_over, C => 
        addr_over, Y => \U1/N_878\);
    
    \U1/cnt_daly_RNO_2[10]\ : NOR3C
      port map(A => \U1/cnt_daly[8]_net_1\, B => 
        \U1/cnt_daly[9]_net_1\, C => \U1/cnt_daly[7]_net_1\, Y
         => \U1/m22_m4_0_a2_3\);
    
    \U0/cnt_rc_n3\ : AX1
      port map(A => \U0/N_130\, B => \U0/cnt_rc_7_0_net_1\, C => 
        \U0/N_59\, Y => \U0/cnt_rc_n3_net_1\);
    
    \U3/data_recive[3]\ : DFN1C0
      port map(D => \U3/data_recive_12[3]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[3]\);
    
    \U3/un7_cnt_1_I_28\ : XOR2
      port map(A => \U3/N_3\, B => \U3/cnt[10]_net_1\, Y => 
        \U3/I_28\);
    
    \U1/ad_once_over\ : DFN1E0C0
      port map(D => \U1/pr_state[4]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1092\, Q => ad_once_over);
    
    \U3/un7_cnt_1_I_18\ : AND3
      port map(A => \U3/cnt[3]_net_1\, B => \U3/cnt[4]_net_1\, C
         => \U3/cnt[5]_net_1\, Y => \U3/DWACT_FINC_E[2]\);
    
    \U5/data_send_RNO_28[4]\ : MX2
      port map(A => \data_all[228]\, B => \data_all[236]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_455\);
    
    \U1/data_all[33]\ : DFN1E0C0
      port map(D => \U1/N_154\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[33]\);
    
    \U1/data_all[142]\ : DFN1E0C0
      port map(D => \U1/N_19\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[142]\);
    
    \U1/cnt_daly_RNIV4081[10]\ : NOR3C
      port map(A => \U1/cnt_daly[9]_net_1\, B => 
        \U1/cnt_daly[10]_net_1\, C => \U1/cnt_daly[7]_net_1\, Y
         => \U1/m20_m6_0_a2_4\);
    
    \U1/data_filter_RNO_1[0]\ : XA1A
      port map(A => \U1/data_filter[0]_net_1\, B => \data_ad[0]\, 
        C => \U1/pr_state_0[5]_net_1\, Y => \U1/N_905\);
    
    \U5/data_send_RNO[4]\ : MX2A
      port map(A => \U5/i67_mux\, B => \U5/N_48_0\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[4]\);
    
    \U3/cnt_RNIOGS11[0]\ : NOR3A
      port map(A => \U3/m27_1\, B => \U3/cnt[3]_net_1\, C => 
        \U3/cnt[0]_net_1\, Y => \U3/m106_7\);
    
    \U1/delay_channel1\ : DFN1E1C0
      port map(D => \U1/pr_state[0]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1838\, Q => 
        \U1/delay_channel1_net_1\);
    
    \U2/cnt[11]\ : DFN1C0
      port map(D => \U2/cnt_n11_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[11]_net_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I80_Y_0\ : AO1
      port map(A => \U1/ADD_14x14_fast_I80_un1_Y_0\, B => 
        \U1/N264\, C => \U1/N263\, Y => 
        \U1/ADD_14x14_fast_I80_Y_0\);
    
    \U1/data_all_RNO_0[224]\ : AO1C
      port map(A => \data_all[224]\, B => \U1/N_837_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_i_0_0_0[224]\);
    
    \U1/data_all_RNO_0[164]\ : AO1C
      port map(A => \data_all[164]\, B => \U1/N_838\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m182_i_0_0\);
    
    \U3/un7_cnt_1_I_23\ : XOR2
      port map(A => \U3/N_5\, B => \U3/cnt[8]_net_1\, Y => 
        \U3/I_23\);
    
    \U3/un7_cnt_1_I_13\ : AND3
      port map(A => \U3/DWACT_FINC_E[0]\, B => \U3/cnt[3]_net_1\, 
        C => \U3/cnt[4]_net_1\, Y => \U3/N_8\);
    
    \U1/data_all[162]\ : DFN1E0C0
      port map(D => \U1/N_1805\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[162]\);
    
    \U2/cnt_25\ : NOR2B
      port map(A => \U2/cnt[11]_net_1\, B => 
        \U2/cnt_0_sqmuxa_net_1\, Y => \U2/N_152\);
    
    \U1/data_filter_RNO_0[6]\ : AO1D
      port map(A => \U1/data_filter[8]_net_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, 
        Y => \U1/m51_0_0_0\);
    
    \U1/data_all_RNO_0[56]\ : AO1C
      port map(A => \data_all[56]\, B => \U1/N_831_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[56]\);
    
    \U1/data_all_RNO_0[153]\ : NOR2A
      port map(A => \U1/N_842\, B => \data_all[153]\, Y => 
        \U1/N_2231\);
    
    \U1/data_all[210]\ : DFN1E0C0
      port map(D => \U1/N_1777\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[210]\);
    
    \U1/data_all[114]\ : DFN1E0C0
      port map(D => \U1/N_368\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[114]\);
    
    \U1/cnt_receive_over_1_sqmuxa\ : NOR2
      port map(A => receive_over, B => addr_over, Y => 
        \U1/cnt_receive_over_1_sqmuxa_net_1\);
    
    \U2/cnt_n5\ : XA1
      port map(A => \U2/cnt[5]_net_1\, B => \U2/cnt_c4_net_1\, C
         => \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n5_net_1\);
    
    \sts_pad/U0/U0\ : IOPAD_IN
      port map(PAD => sts, Y => \sts_pad/U0/NET1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I97_Y\ : XOR3
      port map(A => \U1/data_filter[9]_net_1\, B => \data_ad[9]\, 
        C => \U1/N321\, Y => \U1/un2_data_filter[9]\);
    
    \U1/data_all_RNO_0[59]\ : NOR2A
      port map(A => \U1/N_831\, B => \data_all[59]\, Y => 
        \U1/N_2139\);
    
    \U1/data_all_RNO[65]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[1]_net_1\, 
        C => \U1/m249_i_0_0\, Y => \U1/N_165\);
    
    \U1/data_all_RNO[109]\ : OA1B
      port map(A => \U1/N_829_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/data_all_3_i_0_0_0[109]\, Y => \U1/N_1610\);
    
    \U1/cnt_daly_RNO[0]\ : NOR2
      port map(A => \U1/cnt_daly[0]_net_1\, B => 
        \U1/pr_state[7]_net_1\, Y => \U1/N_42\);
    
    \U1/data_all_RNO[147]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/m109_0_i_0_0\, Y => \U1/N_122\);
    
    \U1/data_all_RNO_0[213]\ : AO1C
      port map(A => \data_all[213]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[213]\);
    
    \U1/cnt_daly_RNI1MV22[8]\ : NOR3C
      port map(A => \U1/cnt_daly[6]_net_1\, B => 
        \U1/cnt_daly[8]_net_1\, C => \U1/m20_m6_0_a2_4\, Y => 
        \U1/m20_m6_0_a2_6\);
    
    \U1/data_all_RNO_0[18]\ : AO1C
      port map(A => \data_all[18]\, B => \U1/N_836_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m159_0_i_0_0\);
    
    \U1/data_all_RNO_0[157]\ : AO1C
      port map(A => \data_all[157]\, B => \U1/N_842\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m79_0_i_i_0\);
    
    \U5/data_send_RNO_4[4]\ : MX2C
      port map(A => \U5/N_495\, B => \U5/N_503\, S => 
        \U5/cnt[2]_net_1\, Y => \U5/N_533\);
    
    \U5/data_send_RNO_26[1]\ : MX2
      port map(A => \data_all[193]\, B => \data_all[201]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_436\);
    
    \U5/data_send[7]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[7]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[7]\);
    
    \U3/data_recive_RNO_0[6]\ : NOR2A
      port map(A => \data_recive[6]\, B => send_over, Y => 
        \U3/m81_0\);
    
    \U2/cnt_n2\ : XA1A
      port map(A => \U2/N_7\, B => \U2/cnt[2]_net_1\, C => 
        \U2/cnt_0_sqmuxa_net_1\, Y => \U2/cnt_n2_net_1\);
    
    \U2/cnt[5]\ : DFN1C0
      port map(D => \U2/cnt_n5_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U2/cnt[5]_net_1\);
    
    \U5/pr_state_RNO_2[0]\ : OR2
      port map(A => send_over, B => \U5/pr_state[1]_net_1\, Y => 
        \U5/N_7\);
    
    \U5/data_send_RNO_2[7]\ : MX2
      port map(A => \U5/N_466\, B => \U5/N_474\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_522\);
    
    \U3/data_recive_RNO_4[5]\ : NOR2A
      port map(A => \U3/cnt[8]_net_1\, B => \U3/cnt[0]_net_1\, Y
         => \U3/m47_1\);
    
    \U1/m206_i_0_o2_0\ : OR2A
      port map(A => \addr_c[0]\, B => \U1/I_5_0\, Y => \U1/N_819\);
    
    \U1/data_all_RNO[48]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[48]\, Y => \U1/N_702\);
    
    \U1/data_all_RNO_1[58]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_831\, 
        Y => \U1/N_2142\);
    
    \U1/m125_0_0_i_o2\ : OR2
      port map(A => \U1/m125_0_0_i_o2_0_net_1\, B => \U1/N_817\, 
        Y => \U1/N_836\);
    
    \U1/data_all_RNO_0[211]\ : NOR2A
      port map(A => \U1/N_840\, B => \data_all[211]\, Y => 
        \U1/N_1029\);
    
    \U1/data_all_RNO_0[11]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[11]\, Y => 
        \U1/N_1075\);
    
    \U1/cnt_daly_RNO[6]\ : XA1C
      port map(A => \U1/cnt_daly[6]_net_1\, B => \U1/N_849\, C
         => \U1/pr_state[7]_net_1\, Y => \U1/N_806\);
    
    \ce_pad/U0/U0\ : IOPAD_TRI
      port map(D => \ce_pad/U0/NET1\, E => \ce_pad/U0/NET2\, PAD
         => ce);
    
    \U1/data_all_RNO_0[73]\ : AO1C
      port map(A => \data_all[73]\, B => \U1/N_833\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m225_i_0_0\);
    
    \U2/cnt_RNI7F1T[11]\ : NOR3C
      port map(A => \U2/cnt[4]_net_1\, B => \U2/cnt[11]_net_1\, C
         => \U2/tx_uart38_10_1\, Y => \U2/tx_uart38_10_3\);
    
    \U1/data_all[94]\ : DFN1E0C0
      port map(D => \U1/data_all_3[94]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[94]\);
    
    \U5/data_send[1]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[1]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[1]\);
    
    \U1/data_all_RNO_1[51]\ : NOR2
      port map(A => \U1/data_filter[3]_net_1\, B => \U1/N_831\, Y
         => \U1/N_2152\);
    
    \U5/data_send_RNO_24[6]\ : MX2
      port map(A => \data_all[166]\, B => \data_all[174]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_425\);
    
    \U2/cnt_RNITBU8Q[8]\ : OR3
      port map(A => \U2/un1_tx_uart27_4_2\, B => 
        \U2/un1_tx_uart27_6\, C => \U2/un1_tx_uart27_5\, Y => 
        \U2/un1_tx_uart27\);
    
    \data_in_pad[9]/U0/U1\ : IOIN_IB
      port map(YIN => \data_in_pad[9]/U0/NET1\, Y => 
        \data_in_c[9]\);
    
    \U1/data_all[90]\ : DFN1E0C0
      port map(D => \U1/N_1775\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[90]\);
    
    \U1/data_all[185]\ : DFN1E0C0
      port map(D => \U1/N_411\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[185]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I69_Y\ : AO1
      port map(A => \U1/N268\, B => \U1/N275\, C => \U1/N267\, Y
         => \U1/N326\);
    
    \U3/un7_cnt_1_I_8\ : AND3
      port map(A => \U3/cnt[0]_net_1\, B => \U3/cnt[1]_net_1\, C
         => \U3/cnt[2]_net_1\, Y => \U3/N_10\);
    
    \U1/pr_state_RNO_0[3]\ : OR3
      port map(A => \U1/N_870\, B => \U1/N_866\, C => \U1/N_869\, 
        Y => \U1/m68_i_i_1\);
    
    \U0/ad_over\ : DFN1E0C0
      port map(D => \U0/pr_state[1]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U0/N_137\, Q => ad_over);
    
    \U1/data_all_RNO_0[7]\ : AO1C
      port map(A => \data_all[7]\, B => \U1/N_835_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[7]\);
    
    \U1/data_all[177]\ : DFN1E0C0
      port map(D => \U1/N_395\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[177]\);
    
    \U4/conver_ris3_RNO\ : INV
      port map(A => \U4/conver_ris2_net_1\, Y => 
        \U4/conver_ris2_i\);
    
    \U1/data_filter_RNO[7]\ : OA1C
      port map(A => \U1/pr_state_0[5]_net_1\, B => 
        \U1/un2_data_filter[7]\, C => \U1/m48_0_0_0\, Y => 
        \U1/N_49_0\);
    
    \U1/data_all_RNO_1[74]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_833\, 
        Y => \U1/N_960\);
    
    \U1/data_all_RNO[237]\ : OA1B
      port map(A => \U1/N_837_0\, B => \U1/data_filter[13]_net_1\, 
        C => \U1/m69_i_0_0\, Y => \U1/N_227\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I93_Y\ : XOR3
      port map(A => \U1/data_filter[5]_net_1\, B => \data_ad[5]\, 
        C => \U1/N332\, Y => \U1/un2_data_filter[5]\);
    
    \U1/m253_i_0_o2\ : OR2
      port map(A => \U1/m253_i_0_o2_0_net_1\, B => \U1/N_817\, Y
         => \U1/N_832\);
    
    \U1/data_all[200]\ : DFN1E0C0
      port map(D => \U1/N_2042\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[200]\);
    
    \U1/data_all[104]\ : DFN1E0C0
      port map(D => \U1/N_50\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[104]\);
    
    \U1/data_all[38]\ : DFN1E0C0
      port map(D => \U1/N_1811\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[38]\);
    
    \rc_pad/U0/U0\ : IOPAD_TRI
      port map(D => \rc_pad/U0/NET1\, E => \rc_pad/U0/NET2\, PAD
         => rc);
    
    \U1/data_all_RNO[58]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2141\, C
         => \U1/N_2142\, Y => \U1/N_686\);
    
    \U3/data_recive[2]\ : DFN1C0
      port map(D => \U3/data_recive_12[2]\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \data_recive[2]\);
    
    \U1/data_all[96]\ : DFN1E0C0
      port map(D => \U1/N_1615\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[96]\);
    
    \U5/data_send_RNO_18[1]\ : MX2
      port map(A => \data_all[65]\, B => \data_all[73]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_372\);
    
    \U1/data_filter[6]\ : DFN1E0C0
      port map(D => \U1/N_52_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[6]_net_1\);
    
    \U1/data_all_RNO[131]\ : OA1B
      port map(A => \U1/N_841_0\, B => \U1/data_filter[3]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[131]\, Y => \U1/N_78\);
    
    \U3/data_recive_RNO_0[7]\ : NOR2A
      port map(A => \data_recive[7]\, B => send_over, Y => 
        \U3/m72_0\);
    
    \U5/data_send_RNO_7[6]\ : MX2
      port map(A => \U5/N_361\, B => \U5/N_369\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_473\);
    
    \U5/data_send_RNO_16[2]\ : MX2
      port map(A => \data_all[34]\, B => \data_all[42]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_357\);
    
    \U5/data_send_RNO[6]\ : MX2A
      port map(A => \U5/i71_mux\, B => \U5/N_34_0\, S => 
        \U5/cnt[4]_net_1\, Y => \U5/un58_data_send[6]\);
    
    \U4/nx_state[1]\ : DLN0P1C1
      port map(D => \GND\, G => \U4/N_24\, PRE => 
        \U4/nx_state_RNO_0[1]_net_1\, CLR => 
        \U4/nx_state_RNO[1]_net_1\, Q => \U4/nx_state[1]_net_1\);
    
    \U2/cnt_RNI8PAD2[4]\ : NOR3C
      port map(A => \U2/tx_uart36_7\, B => \U2/tx_uart36_6\, C
         => \U2/tx_uart36_8\, Y => \U2/tx_uart36\);
    
    \U1/cnt_daly_RNO_0[10]\ : NOR3B
      port map(A => \U1/m22_m4_0_a2_4\, B => \U1/m22_m4_0_a2_3\, 
        C => \U1/N_846\, Y => \U1/m22_N_11_mux\);
    
    \U2/cnt_n0\ : NOR2A
      port map(A => \U2/cnt_0_sqmuxa_net_1\, B => 
        \U2/cnt[0]_net_1\, Y => \U2/cnt_n0_net_1\);
    
    \U0/pr_state[0]\ : DFN1C0
      port map(D => \U0/pr_state_RNO_0[0]_net_1\, CLK => 
        sys_clk_c, CLR => sys_rest_c, Q => \U0/pr_state[0]_net_1\);
    
    \sys_clk_pad/U0/U0\ : IOPAD_IN
      port map(PAD => sys_clk, Y => \sys_clk_pad/U0/NET1\);
    
    \U1/data_all_RNO_0[236]\ : NOR2A
      port map(A => \U1/N_837\, B => \data_all[236]\, Y => 
        \U1/N_983\);
    
    \U1/data_all_RNO[233]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_911\, C
         => \U1/N_912\, Y => \U1/N_223\);
    
    \U1/cnt_daly_RNO[8]\ : NOR3A
      port map(A => \U1/N_852\, B => \U1/pr_state[7]_net_1\, C
         => \U1/N_2303\, Y => \U1/N_810\);
    
    \U5/data_send[2]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[2]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[2]\);
    
    \U4/conver_ris_RNO\ : NOR2B
      port map(A => \U4/conver_ris3_i_0\, B => 
        \U4/conver_ris2_net_1\, Y => \U4/conver_ris_2\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I52_Y\ : AO1
      port map(A => \U1/N248\, B => \U1/N245\, C => \U1/N244\, Y
         => \U1/N271\);
    
    \U0/pr_state_RNIF752[5]\ : AO1A
      port map(A => addr_over, B => \U0/pr_state[5]_net_1\, C => 
        \U0/N_137\, Y => \U0/un1_pr_state_5\);
    
    \U1/data_all_3_i_0_0_o2[126]\ : OR3
      port map(A => \U1/N_818\, B => \U1/N_820\, C => 
        \addr_c_0[0]\, Y => \U1/N_830\);
    
    \U5/data_send_RNO_15[0]\ : MX2
      port map(A => \data_all[16]\, B => \data_all[24]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_347\);
    
    \U1/data_all[95]\ : DFN1E0C0
      port map(D => \U1/data_all_3[95]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[95]\);
    
    \U1/data_all[195]\ : DFN1E0C0
      port map(D => \U1/N_201\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[195]\);
    
    \U1/data_all_RNO[191]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \data_all[191]\, 
        C => \U1/N_844_0\, Y => \U1/N_51\);
    
    \U1/data_all_RNO[94]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_834_0\, C
         => \data_all[94]\, Y => \U1/data_all_3[94]\);
    
    \U5/data_send_RNO_12[6]\ : MX2
      port map(A => \U5/N_441\, B => \U5/N_449\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_513\);
    
    \U1/pr_state_RNI281B1[6]\ : OR3
      port map(A => \U1/pr_state[2]_net_1\, B => 
        \U1/pr_state[0]_net_1\, C => \U1/pr_state[6]_net_1\, Y
         => \U1/N_857\);
    
    \U1/data_all_RNO_0[74]\ : NOR2A
      port map(A => \U1/N_833\, B => \data_all[74]\, Y => 
        \U1/N_959\);
    
    \U1/data_all_RNO_0[212]\ : AO1C
      port map(A => \data_all[212]\, B => \U1/N_840_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[212]\);
    
    \U1/data_filter_RNO_0[8]\ : AO1D
      port map(A => \U1/data_filter[10]_net_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/pr_state_0[7]_net_1\, 
        Y => \U1/data_filter_4_i_0_0_0[8]\);
    
    \U5/data_send_RNO_19[2]\ : MX2
      port map(A => \data_all[82]\, B => \data_all[90]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_381\);
    
    \U4/addr_RNO[3]\ : XA1
      port map(A => \addr_c[3]\, B => \U4/N_9_0\, C => 
        \U4/pr_state[0]_net_1\, Y => \U4/addr_n3\);
    
    \U3/un7_cnt_1_I_26\ : AX1C
      port map(A => \U3/cnt[8]_net_1\, B => \U3/DWACT_FINC_E[4]\, 
        C => \U3/cnt[9]_net_1\, Y => \U3/I_26\);
    
    \U5/data_send_RNO_17[3]\ : MX2
      port map(A => \data_all[51]\, B => \data_all[59]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_366\);
    
    \U3/un7_cnt_1_I_16\ : AND3
      port map(A => \U3/DWACT_FINC_E[0]\, B => 
        \U3/DWACT_FINC_E[1]\, C => \U3/cnt[5]_net_1\, Y => 
        \U3/N_7\);
    
    \U3/data_recive_RNO_1[7]\ : NOR3C
      port map(A => \U3/m22_2\, B => \U3/m22_1\, C => 
        \U3/N_125_mux\, Y => \U3/data_recive30\);
    
    \U2/tx_uart_RNO_6\ : NOR2B
      port map(A => \U2/parity_check_8_sqmuxa\, B => 
        \data_send[7]\, Y => \U2/data_send_m[7]\);
    
    \U1/delay_channel1_RNO_0\ : NOR2B
      port map(A => \U1/pr_state[0]_net_1\, B => \addr_c[0]\, Y
         => \U1/m101_i_0_a3_0_0\);
    
    \U3/data_recive_RNO_2[2]\ : NOR3B
      port map(A => \U3/cnt[0]_net_1\, B => \U3/m27_1\, C => 
        \U3/cnt[3]_net_1\, Y => \U3/m70_5\);
    
    \U1/data_all[32]\ : DFN1E0C0
      port map(D => \U1/N_1806\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[32]\);
    
    \U0/data_ad[10]\ : DFN1E0C0
      port map(D => \U0/data_ad_4[10]\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U0/un1_pr_state_5\, Q => \data_ad[10]\);
    
    \U5/vld_send_RNO\ : NOR2A
      port map(A => \U5/pr_state[1]_net_1\, B => \U5/N_138_mux\, 
        Y => \U5/N_78\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I0_CO1\ : NOR2B
      port map(A => \data_ad[0]\, B => \U1/data_filter[0]_net_1\, 
        Y => \U1/N176\);
    
    \U1/data_all_RNO_0[133]\ : AO1C
      port map(A => \data_all[133]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[133]\);
    
    \U1/data_all_RNO[219]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1017\, C
         => \U1/N_1018\, Y => \U1/N_170\);
    
    \U0/pr_state_RNI0EH[1]\ : NOR2
      port map(A => \U0/pr_state[1]_net_1\, B => 
        \U0/pr_state[5]_net_1\, Y => \U0/N_137\);
    
    \U5/data_send_RNO_21[0]\ : MX2
      port map(A => \data_all[112]\, B => \data_all[120]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_395\);
    
    \U1/receive_on_RNIOEGQ\ : OR2B
      port map(A => receive_on, B => \U1/pr_state[7]_net_1\, Y
         => \U1/N_860\);
    
    \U2/send_RNO\ : OR2B
      port map(A => \U2/idle_send_net_1\, B => vld_send, Y => 
        \U2/un5_vld_send\);
    
    \U2/cnt_RNIH1K9_1[9]\ : NOR2
      port map(A => \U2/cnt[9]_net_1\, B => \U2/cnt[4]_net_1\, Y
         => \U2/N_176\);
    
    \U1/data_all[214]\ : DFN1E0C0
      port map(D => \U1/N_182\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[214]\);
    
    \U0/conver_ris2\ : DFN1C0
      port map(D => \U0/conver_ris1_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, Q => \U0/conver_ris2_net_1\);
    
    \U5/data_send_RNO_6[0]\ : MX2
      port map(A => \U5/N_339\, B => \U5/N_347\, S => 
        \U5/cnt[1]_net_1\, Y => \U5/N_459\);
    
    \U5/data_send_RNO_0[7]\ : MX2A
      port map(A => \U5/N_522\, B => \U5/N_538\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/i58_mux\);
    
    \U5/data_send[4]\ : DFN1E1C0
      port map(D => \U5/un58_data_send[4]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U5/pr_state[0]_net_1\, Q => 
        \data_send[4]\);
    
    \U1/data_all_RNO[5]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1086\, C
         => \U1/N_1087\, Y => \U1/N_253\);
    
    \U1/data_all_RNO_0[137]\ : AO1C
      port map(A => \data_all[137]\, B => \U1/N_841\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[137]\);
    
    \U1/data_all_RNO[79]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_833\, C
         => \data_all[79]\, Y => \U1/data_all_3[79]\);
    
    \U1/data_all_RNO_0[82]\ : NOR2A
      port map(A => \U1/N_834\, B => \data_all[82]\, Y => 
        \U1/N_1047\);
    
    \U5/data_send_RNO_18[2]\ : MX2
      port map(A => \data_all[66]\, B => \data_all[74]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_373\);
    
    \U2/tx_uart_RNO_8\ : AO1
      port map(A => \U2/parity_check_5_sqmuxa\, B => 
        \data_send[4]\, C => \U2/data_send_m[6]\, Y => 
        \U2/tx_uart_11_iv_3\);
    
    \U1/cnt_daly[8]\ : DFN1E0C0
      port map(D => \U1/N_810\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1090\, Q => \U1/cnt_daly[8]_net_1\);
    
    \U4/conver_ris_RNIK7T62\ : MX2B
      port map(A => \U4/N_22\, B => \U4/N_10_0\, S => 
        ad_once_over, Y => \U4/N_23\);
    
    \U4/pr_state_RNIMCFF2[1]\ : NOR2
      port map(A => \U4/N_23\, B => \U4/pr_state[1]_net_1\, Y => 
        \U4/N_24\);
    
    \U2/cnt_RNISS7J[9]\ : NOR2B
      port map(A => \U2/N_164\, B => \U2/N_163\, Y => \U2/N_180\);
    
    \U1/data_all[141]\ : DFN1E0C0
      port map(D => \U1/N_97\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[141]\);
    
    \U3/cnt_RNIJFUG[5]\ : NOR2A
      port map(A => \U3/cnt[8]_net_1\, B => \U3/cnt[5]_net_1\, Y
         => \U3/m36_1\);
    
    \U1/data_all_RNO_1[10]\ : NOR2
      port map(A => \U1/data_filter[10]_net_1\, B => \U1/N_835\, 
        Y => \U1/N_2296\);
    
    \U1/data_all[238]\ : DFN1E0C0
      port map(D => \U1/N_160\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[238]\);
    
    \U1/data_all_RNO[114]\ : OA1B
      port map(A => \U1/N_830_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[114]\, Y => \U1/N_368\);
    
    \U1/data_all_RNO[211]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1029\, C
         => \U1/N_1030\, Y => \U1/N_192\);
    
    \U5/data_send_RNO_20[6]\ : MX2
      port map(A => \data_all[102]\, B => \data_all[110]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_393\);
    
    \U2/cnt_RNI1J3G1[0]\ : NOR2B
      port map(A => \U2/tx_uart35_0_a2_0_1\, B => \U2/N_172\, Y
         => \U2/N_192\);
    
    \U1/data_all_RNO[162]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/m71_i_0_0\, Y => \U1/N_1805\);
    
    \U1/data_all[161]\ : DFN1E0C0
      port map(D => \U1/N_1815\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[161]\);
    
    \addr_pad[1]/U0/U1\ : IOTRI_OB_EB
      port map(D => \addr_c[1]\, E => \VCC\, DOUT => 
        \addr_pad[1]/U0/NET1\, EOUT => \addr_pad[1]/U0/NET2\);
    
    \U5/pr_state[1]\ : DFN1C0
      port map(D => \U5/pr_state_RNO[1]_net_1\, CLK => sys_clk_c, 
        CLR => sys_rest_c, Q => \U5/pr_state[1]_net_1\);
    
    \U1/data_filter_RNO[10]\ : OA1C
      port map(A => \U1/pr_state_0[5]_net_1\, B => 
        \U1/un2_data_filter[10]\, C => 
        \U1/data_filter_4_i_0_0_0[10]\, Y => \U1/N_37\);
    
    \U1/data_all_RNO[89]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2133\, C
         => \U1/N_2134\, Y => \U1/N_360\);
    
    \U5/data_send_RNO_1[2]\ : MX2A
      port map(A => \U5/N_535\, B => \U5/N_61_0\, S => 
        \U5/cnt[3]_net_1\, Y => \U5/N_62_0\);
    
    \U1/data_all[31]\ : DFN1E0C0
      port map(D => \U1/data_all_3[31]\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1091\, Q => \data_all[31]\);
    
    \U1/data_all_RNO[210]\ : OA1B
      port map(A => \U1/N_840_0\, B => \U1/data_filter[2]_net_1\, 
        C => \U1/data_all_3_0_i_0_0[210]\, Y => \U1/N_1777\);
    
    \U1/data_all[37]\ : DFN1E0C0
      port map(D => \U1/N_1810\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[37]\);
    
    \rx_uart_pad/U0/U1\ : IOIN_IB
      port map(YIN => \rx_uart_pad/U0/NET1\, Y => rx_uart_c);
    
    \U1/pr_state_RNISSL91[7]\ : OR2
      port map(A => \U1/N_119\, B => \U1/pr_state[7]_net_1\, Y
         => \U1/N_793\);
    
    \U1/delay_channel1_RNI00551\ : OR2A
      port map(A => \U4.N_31\, B => \U1/delay_channel1_net_1\, Y
         => \U1/N_856\);
    
    \U1/data_filter_RNO[2]\ : OA1C
      port map(A => \U1/pr_state[5]_net_1\, B => 
        \U1/un2_data_filter[2]\, C => 
        \U1/data_filter_4_i_0_0_0[2]\, Y => \U1/N_45\);
    
    \U1/data_all[8]\ : DFN1E0C0
      port map(D => \U1/N_246\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[8]\);
    
    \U1/data_filter_RNO_0[0]\ : NOR2
      port map(A => \U1/data_filter[2]_net_1\, B => 
        \U1/pr_state[5]_net_1\, Y => \U1/N_906\);
    
    \U1/data_all_RNO_1[235]\ : NOR2
      port map(A => \U1/data_filter[11]_net_1\, B => \U1/N_837_0\, 
        Y => \U1/N_910\);
    
    \U3/data_recive_RNO[5]\ : MX2
      port map(A => \U3/m83_0\, B => rx_uart_c, S => 
        \U3/data_recive28\, Y => \U3/data_recive_12[5]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I26_Y\ : MAJ3
      port map(A => \U1/N188\, B => \U1/data_filter[5]_net_1\, C
         => \data_ad[5]\, Y => \U1/N242\);
    
    \U1/data_all_RNO_0[0]\ : AO1C
      port map(A => \data_all[0]\, B => \U1/N_835_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_0_i_0[0]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I77_un1_Y_0\ : NOR3C
      port map(A => \U1/N243\, B => \U1/N239\, C => \U1/N258\, Y
         => \U1/ADD_14x14_fast_I77_un1_Y_0\);
    
    \U1/data_all_RNO_0[161]\ : AO1C
      port map(A => \data_all[161]\, B => \U1/N_838_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m188_i_0_0\);
    
    \U3/data_recive_RNO_0[4]\ : NOR2A
      port map(A => \data_recive[4]\, B => send_over, Y => 
        \U3/m85_0\);
    
    \U1/pr_state_RNO_0[6]\ : AO1
      port map(A => \U1/N_1084\, B => \U1/pr_state_0[5]_net_1\, C
         => \U1/N_878\, Y => \U1/m77_i_0_0\);
    
    \U3/cnt_4[3]\ : XA1
      port map(A => \U3/N_10\, B => \U3/cnt[3]_net_1\, C => 
        \U3/recive_net_1\, Y => \U3/cnt_4[3]_net_1\);
    
    \U1/data_all_RNO[144]\ : OA1B
      port map(A => \U1/N_842_0\, B => \U1/data_filter[0]_net_1\, 
        C => \U1/m118_0_i_1_0\, Y => \U1/N_1794\);
    
    \U1/data_all[23]\ : DFN1E0C0
      port map(D => \U1/N_1788\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[23]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I17_Y\ : NOR2B
      port map(A => \U1/N207\, B => \U1/N204\, Y => \U1/N233\);
    
    \U1/data_all[204]\ : DFN1E0C0
      port map(D => \U1/N_100\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[204]\);
    
    \U1/data_all_RNO[172]\ : OA1B
      port map(A => \U1/N_838_0\, B => \U1/data_filter[12]_net_1\, 
        C => \U1/m156_i_0_0\, Y => \U1/N_331\);
    
    \U1/data_all[228]\ : DFN1E0C0
      port map(D => \U1/N_215\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[228]\);
    
    \U1/cnt_daly_RNIP7VQ[2]\ : NOR2B
      port map(A => \U1/cnt_daly[2]_net_1\, B => 
        \U1/cnt_daly[3]_net_1\, Y => \U1/m20_m6_0_a2_1\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I22_Y\ : MAJ3
      port map(A => \U1/N194\, B => \U1/data_filter[7]_net_1\, C
         => \data_ad[7]\, Y => \U1/N238\);
    
    \U1/data_all_3_i_0_0_o2_0[126]\ : OR3
      port map(A => \U1/N_818\, B => \U1/N_820\, C => 
        \addr_c_0[0]\, Y => \U1/N_830_0\);
    
    \U1/vld_whole\ : DFN1E0C0
      port map(D => \U1/N_858\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1093\, Q => vld_whole);
    
    \U1/conver\ : DFN1E0C0
      port map(D => \U1/pr_state[6]_net_1\, CLK => sys_clk_c, CLR
         => sys_rest_c, E => \U1/N_1095\, Q => conver_top);
    
    \U1/data_all_RNO[43]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2197\, C
         => \U1/N_2198\, Y => \U1/N_284\);
    
    \U3/cnt_RNIS0VF_0[10]\ : NOR2A
      port map(A => \U3/cnt[5]_net_1\, B => \U3/cnt[10]_net_1\, Y
         => \U3/m11_3\);
    
    \U1/data_all_RNO_0[10]\ : NOR2A
      port map(A => \U1/N_835\, B => \data_all[10]\, Y => 
        \U1/N_2295\);
    
    \U1/data_all[182]\ : DFN1E0C0
      port map(D => \U1/N_405\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[182]\);
    
    \U1/data_all_RNO[152]\ : OA1B
      port map(A => \U1/N_842\, B => \U1/data_filter[8]_net_1\, C
         => \U1/m92_1_i_0_0\, Y => \U1/N_1798\);
    
    \U5/data_send_RNO_22[7]\ : MX2
      port map(A => \data_all[135]\, B => \data_all[143]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_410\);
    
    \U1/data_all_RNO[69]\ : OA1B
      port map(A => \U1/N_833_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/m237_i_0_0\, Y => \U1/N_173\);
    
    \addr_pad[0]/U0/U1\ : IOTRI_OB_EB
      port map(D => \addr_c[0]\, E => \VCC\, DOUT => 
        \addr_pad[0]/U0/NET1\, EOUT => \addr_pad[0]/U0/NET2\);
    
    \U3/rx_fall1\ : DFN1C0
      port map(D => \U3/rx_fall_net_1\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/rx_fall1_net_1\);
    
    \U1/data_filter[2]\ : DFN1E0C0
      port map(D => \U1/N_45\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[2]_net_1\);
    
    \U1/data_all_RNO[186]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2081\, C
         => \U1/N_2082\, Y => \U1/N_413\);
    
    \U5/data_send_RNO_27[2]\ : MX2
      port map(A => \data_all[210]\, B => \data_all[218]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_445\);
    
    \U1/data_all_RNO[3]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_1096\, C
         => \U1/N_1097\, Y => \U1/N_258\);
    
    \U1/pr_state_RNIV2MS[1]\ : NOR2
      port map(A => \U1/pr_state[1]_net_1\, B => 
        \U1/pr_state[2]_net_1\, Y => 
        \U1/pr_state_RNIV2MS[1]_net_1\);
    
    \U1/data_all[9]\ : DFN1E0C0
      port map(D => \U1/N_243\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[9]\);
    
    \U1/data_all_RNO_1[50]\ : NOR2
      port map(A => \U1/data_filter[2]_net_1\, B => \U1/N_831\, Y
         => \U1/N_2154\);
    
    \U3/data_recive_RNO_1[2]\ : NOR3C
      port map(A => \U3/m70_5\, B => \U3/m70_4\, C => \U3/N_29\, 
        Y => \U3/data_recive25\);
    
    \U1/pr_state_0_RNIAOTO2[5]\ : NOR3A
      port map(A => \U1/m85_i_0_a3_1\, B => 
        \U1/pr_state_0[5]_net_1\, C => \U1/N_857\, Y => 
        \U1/N_871\);
    
    \U1/data_filter[5]\ : DFN1E0C0
      port map(D => \U1/N_55_0\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1094\, Q => 
        \U1/data_filter[5]_net_1\);
    
    \U1/data_all[173]\ : DFN1E0C0
      port map(D => \U1/N_333\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[173]\);
    
    \U1/data_all[135]\ : DFN1E0C0
      port map(D => \U1/N_105\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[135]\);
    
    \U1/un14_data_all_I_5\ : XNOR2
      port map(A => \addr_c[0]\, B => \addr_c[1]\, Y => 
        \U1/I_5_0\);
    
    \U1/data_all_RNO_1[82]\ : NOR2
      port map(A => \U1/data_filter[2]_net_1\, B => \U1/N_834\, Y
         => \U1/N_1048\);
    
    \U3/data_recive_RNO_0[3]\ : NOR2A
      port map(A => \data_recive[3]\, B => send_over, Y => 
        \U3/m87_0\);
    
    \U5/data_send_RNO_14[4]\ : MX2
      port map(A => \data_all[4]\, B => \data_all[12]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_343\);
    
    \U1/data_all_RNO[14]\ : NOR3C
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_835_0\, C
         => \data_all[14]\, Y => \U1/data_all_3[14]\);
    
    \U1/data_all_3_0_0_i_o2[92]\ : OR2
      port map(A => \U1/N_826\, B => \U1/N_821\, Y => \U1/N_834\);
    
    \U5/data_send_RNO_27[1]\ : MX2
      port map(A => \data_all[209]\, B => \data_all[217]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_444\);
    
    \U2/cnt_c8\ : NOR2B
      port map(A => \U2/cnt_c7_net_1\, B => \U2/cnt[8]_net_1\, Y
         => \U2/cnt_c8_net_1\);
    
    \U1/data_all_RNO_0[114]\ : AO1C
      port map(A => \data_all[114]\, B => \U1/N_830\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/data_all_3_0_i_0_0[114]\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I91_Y\ : XOR3
      port map(A => \U1/data_filter[3]_net_1\, B => \data_ad[3]\, 
        C => \U1/N275\, Y => \U1/un2_data_filter[3]\);
    
    \U5/data_send_RNO_16[3]\ : MX2
      port map(A => \data_all[35]\, B => \data_all[43]\, S => 
        \U5/cnt[0]_net_1\, Y => \U5/N_358\);
    
    \U3/data_recive_RNO_2[5]\ : NOR3B
      port map(A => \U3/cnt[10]_net_1\, B => \U3/m47_1\, C => 
        \U3/cnt[5]_net_1\, Y => \U3/m47_3\);
    
    \U2/cnt_c1_i_RNIA2GG1\ : NOR2B
      port map(A => \U2/tx_uart38_10_4\, B => \U2/tx_uart38_10_3\, 
        Y => \U2/tx_uart38_10\);
    
    \U1/data_all[99]\ : DFN1E0C0
      port map(D => \U1/N_60\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[99]\);
    
    \U3/cnt[8]\ : DFN1C0
      port map(D => \U3/I_23\, CLK => sys_clk_c, CLR => 
        sys_rest_c, Q => \U3/cnt[8]_net_1\);
    
    \U1/data_all_RNO[76]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_955\, C
         => \U1/N_956\, Y => \U1/N_187\);
    
    \U1/data_all_RNO_1[236]\ : NOR2
      port map(A => \U1/data_filter[12]_net_1\, B => \U1/N_837\, 
        Y => \U1/N_984\);
    
    \U1/data_all_RNO_0[193]\ : AO1C
      port map(A => \data_all[193]\, B => \U1/N_839_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m142_0_i_0\);
    
    \U1/data_all_RNO[28]\ : NOR3A
      port map(A => \U1/pr_state[2]_net_1\, B => \U1/N_2253\, C
         => \U1/N_2254\, Y => \U1/N_765\);
    
    \U0/pr_state_RNO[2]\ : NOR2A
      port map(A => \U0/pr_state[3]_net_1\, B => \U0/sts_ris_i_0\, 
        Y => \U0/pr_state_RNO[2]_net_1\);
    
    \U1/cnt_daly_RNI83HF2[11]\ : NOR3C
      port map(A => \U1/m61_0_i_a3_1_1\, B => \U1/m61_0_i_a3_1_0\, 
        C => \U1/m61_0_i_a3_1_5\, Y => \U1/m61_0_i_a3_1_9\);
    
    \U1/un2_data_filter_ADD_14x14_fast_I13_Y\ : OA1
      port map(A => \U1/data_filter[11]_net_1\, B => 
        \data_ad[11]\, C => \U1/data_filter[12]_net_1\, Y => 
        \U1/N229\);
    
    \U1/data_all_RNO[53]\ : OA1B
      port map(A => \U1/N_831_0\, B => \U1/data_filter[5]_net_1\, 
        C => \U1/data_all_3_0_0_i_0[53]\, Y => \U1/N_48\);
    
    \U1/data_all[192]\ : DFN1E0C0
      port map(D => \U1/N_197\, CLK => sys_clk_c, CLR => 
        sys_rest_c, E => \U1/N_1091\, Q => \data_all[192]\);
    
    \U5/data_send_RNO_5[3]\ : MX2
      port map(A => \U5/N_510\, B => \U5/N_53_0\, S => 
        \U5/cnt_0[2]_net_1\, Y => \U5/N_54_0\);
    
    \U3/rx_down_RNO\ : NOR2A
      port map(A => \U3/rx_fall2_net_1\, B => \U3/rx_fall1_net_1\, 
        Y => \U3/rx_down_1\);
    
    \U1/data_all_3_i_0_0_o2_0[111]\ : OR3A
      port map(A => \addr_c_0[0]\, B => \U1/N_818\, C => 
        \U1/N_820\, Y => \U1/N_829_0\);
    
    \U1/data_all_RNO_0[197]\ : AO1C
      port map(A => \data_all[197]\, B => \U1/N_839_0\, C => 
        \U1/pr_state[2]_net_1\, Y => \U1/m130_0_i_0\);
    
    GND_power_inst1 : GND
      port map( Y => GND_power_net1);

    VCC_power_inst1 : VCC
      port map( Y => VCC_power_net1);


end DEF_ARCH; 
